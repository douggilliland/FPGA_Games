module BLUETOOTH(
	input clk,
	input reg [10:0]din,
	input enable, 
        input RW,
	input Rx,
	output Tx,
	output [10:0]dout,
	output done, 
	output busy,
);

	r
