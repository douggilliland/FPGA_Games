library IEEE;
use IEEE.STD_LOGIC_1164.all;



entity objects_draw is
port 	(
		--////////////////////	Clock Input	 	////////////////////	
	   CLK  					: in std_logic;
		RESETn				: in std_logic;
		oCoord_X				: in integer;
		oCoord_Y				: in integer;
		fell_to_pit			: in std_logic ;
		game_started 		: in std_logic ;
		space_was_pressed : in std_logic ;
		game_over			: in std_logic ;
		bounce_type 		: out std_logic_vector(4 downto 0) ;
		drawing_request	: out std_logic ;
		mVGA_RGB 			: out std_logic_vector(7 downto 0) 
	);
end entity;

architecture behav of objects_draw is 

	-- posting the title
	signal sigSpaceWasPressed : std_logic := '0';
	signal sigGameOver : std_logic := '0';
	-- /posting the title
	--All Purpose :
	signal sig_draw_req : std_logic := '0';
	signal sig_draw_data: std_logic_vector (7 downto 0);
	signal sig_bounce_type : std_logic_vector (4 downto 0);
	
	--signal game_started : std_logic := '0';
	constant game_started_X_bound : integer := 560;
	
	--signal fell_to_pit : std_logic := '0';
	constant fell_to_pit_right_X_bound : integer := 378;
	constant fell_to_pit_left_X_bound : integer := 192;
	constant fell_to_pit_upper_Y_bound : integer := 382;

	constant no_bounce			 		: std_logic_vector (4 downto 0) := "00000";
	constant horizontal_floor 			: std_logic_vector (4 downto 0) := "00001";
	constant left_down_slope 			: std_logic_vector (4 downto 0) := "00010";
	constant left_vertical_wall 		: std_logic_vector (4 downto 0) := "00011";
	constant left_up_slope 				: std_logic_vector (4 downto 0) := "00100";
	constant horizontal_ceiling 		: std_logic_vector (4 downto 0) := "00101";
	constant right_up_slope 			: std_logic_vector (4 downto 0) := "00110";
	constant right_vertical_wall 		: std_logic_vector (4 downto 0) := "00111";
	constant right_down_slope 			: std_logic_vector (4 downto 0) := "01000";
	constant death				 		: std_logic_vector (4 downto 0) := "01001";

	--floor:
	constant floor_start_x 	: integer := 0;
	constant floor_start_y 	: integer := 450;
	constant floor_X_size 	: integer := 640;
	constant floor_Y_size 	: integer := 30;
	constant floor_color  	: std_logic_vector(7 downto 0) := x"e1";
	constant floor_bounce_type : std_logic_vector(4 downto 0) := horizontal_floor;
	signal floor_end_x : integer;
	signal floor_end_y : integer;
	signal floor_drawing_X : std_logic := '0';
	signal floor_drawing_Y : std_logic := '0';
	signal floor_drawing_req : std_logic := '0';
	--/floor
	
	--right_wall:
	constant right_wall_start_x 	: integer := 610;
	constant right_wall_start_y 	: integer := 30;
	constant right_wall_X_size 	: integer := 30;
	constant right_wall_Y_size 	: integer := 420;
	constant right_wall_color  	: std_logic_vector(7 downto 0) := x"d0";
	constant right_wall_bounce_type : std_logic_vector(4 downto 0) := right_vertical_wall;
	signal right_wall_end_x : integer;
	signal right_wall_end_y : integer;
	signal right_wall_drawing_X : std_logic := '0';
	signal right_wall_drawing_Y : std_logic := '0';
	signal right_wall_drawing_req : std_logic := '0';
	--/right_wall
	
	--left_wall:
	constant left_wall_start_x 	: integer := 0;
	constant left_wall_start_y 	: integer := 30;
	constant left_wall_X_size 	: integer := 30;
	constant left_wall_Y_size 	: integer := 420;
	constant left_wall_color  	: std_logic_vector(7 downto 0) := x"d0";
	constant left_wall_bounce_type : std_logic_vector(4 downto 0) := left_vertical_wall;
	signal left_wall_end_x : integer;
	signal left_wall_end_y : integer;
	signal left_wall_drawing_X : std_logic := '0';
	signal left_wall_drawing_Y : std_logic := '0';
	signal left_wall_drawing_req : std_logic := '0';
	--/left_wall
	
	--ceiling:
	constant ceiling_start_x 	: integer := 0;
	constant ceiling_start_y 	: integer := 0;
	constant ceiling_X_size 	: integer := 640;
	constant ceiling_Y_size 	: integer := 30;
	constant ceiling_color  	: std_logic_vector(7 downto 0) := x"d0";
	constant ceiling_bounce_type : std_logic_vector(4 downto 0) := horizontal_ceiling;
	signal ceiling_end_x : integer;
	signal ceiling_end_y : integer;
	signal ceiling_drawing_X : std_logic := '0';
	signal ceiling_drawing_Y : std_logic := '0';
	signal ceiling_drawing_req : std_logic := '0';
	--/ceiling
	
	--left_down_slope:
	constant left_down_slope_start_x 	: integer := 30;
	constant left_down_slope_start_y 	: integer := 310;
	constant left_down_slope_X_size 	: integer := 70;
	constant left_down_slope_Y_size 	: integer := 70;
	constant left_down_slope_color  	: std_logic_vector(7 downto 0) := x"83";
	constant left_down_slope_bounce_type : std_logic_vector(4 downto 0) := left_down_slope;
	signal left_down_slope_end_x : integer;
	signal left_down_slope_end_y : integer;
	signal left_down_slope_drawing_X : std_logic := '0';
	signal left_down_slope_drawing_Y : std_logic := '0';
	signal left_down_slope_drawing_req : std_logic := '0';
	signal left_down_slope_Coord_X : integer := 0;-- offset from start position 
	signal left_down_slope_Coord_Y : integer := 0;
	--/left_down_slope
	
	type left_down_slope_object_form is array (0 to left_down_slope_Y_size - 1 , 0 to left_down_slope_X_size - 1) of std_logic;
	constant left_down_slope_object : left_down_slope_object_form := (
("1000000000000000000000000000000000000000000000000000000000000000000000"),
("1100000000000000000000000000000000000000000000000000000000000000000000"),
("1110000000000000000000000000000000000000000000000000000000000000000000"),
("1111000000000000000000000000000000000000000000000000000000000000000000"),
("1111100000000000000000000000000000000000000000000000000000000000000000"),
("1111110000000000000000000000000000000000000000000000000000000000000000"),
("1111111000000000000000000000000000000000000000000000000000000000000000"),
("1111111100000000000000000000000000000000000000000000000000000000000000"),
("1111111110000000000000000000000000000000000000000000000000000000000000"),
("1111111111000000000000000000000000000000000000000000000000000000000000"),
("1111111111100000000000000000000000000000000000000000000000000000000000"),
("1111111111110000000000000000000000000000000000000000000000000000000000"),
("1111111111111000000000000000000000000000000000000000000000000000000000"),
("1111111111111100000000000000000000000000000000000000000000000000000000"),
("1111111111111110000000000000000000000000000000000000000000000000000000"),
("1111111111111111000000000000000000000000000000000000000000000000000000"),
("1111111111111111100000000000000000000000000000000000000000000000000000"),
("1111111111111111110000000000000000000000000000000000000000000000000000"),
("1111111111111111111000000000000000000000000000000000000000000000000000"),
("1111111111111111111100000000000000000000000000000000000000000000000000"),
("1111111111111111111110000000000000000000000000000000000000000000000000"),
("1111111111111111111111000000000000000000000000000000000000000000000000"),
("1111111111111111111111100000000000000000000000000000000000000000000000"),
("1111111111111111111111110000000000000000000000000000000000000000000000"),
("1111111111111111111111111000000000000000000000000000000000000000000000"),
("1111111111111111111111111100000000000000000000000000000000000000000000"),
("1111111111111111111111111110000000000000000000000000000000000000000000"),
("1111111111111111111111111111000000000000000000000000000000000000000000"),
("1111111111111111111111111111100000000000000000000000000000000000000000"),
("1111111111111111111111111111110000000000000000000000000000000000000000"),
("1111111111111111111111111111111000000000000000000000000000000000000000"),
("1111111111111111111111111111111100000000000000000000000000000000000000"),
("1111111111111111111111111111111110000000000000000000000000000000000000"),
("1111111111111111111111111111111111000000000000000000000000000000000000"),
("1111111111111111111111111111111111100000000000000000000000000000000000"),
("1111111111111111111111111111111111110000000000000000000000000000000000"),
("1111111111111111111111111111111111111000000000000000000000000000000000"),
("1111111111111111111111111111111111111100000000000000000000000000000000"),
("1111111111111111111111111111111111111110000000000000000000000000000000"),
("1111111111111111111111111111111111111111000000000000000000000000000000"),
("1111111111111111111111111111111111111111100000000000000000000000000000"),
("1111111111111111111111111111111111111111110000000000000000000000000000"),
("1111111111111111111111111111111111111111111000000000000000000000000000"),
("1111111111111111111111111111111111111111111100000000000000000000000000"),
("1111111111111111111111111111111111111111111110000000000000000000000000"),
("1111111111111111111111111111111111111111111111000000000000000000000000"),
("1111111111111111111111111111111111111111111111100000000000000000000000"),
("1111111111111111111111111111111111111111111111110000000000000000000000"),
("1111111111111111111111111111111111111111111111111000000000000000000000"),
("1111111111111111111111111111111111111111111111111100000000000000000000"),
("1111111111111111111111111111111111111111111111111110000000000000000000"),
("1111111111111111111111111111111111111111111111111111000000000000000000"),
("1111111111111111111111111111111111111111111111111111100000000000000000"),
("1111111111111111111111111111111111111111111111111111110000000000000000"),
("1111111111111111111111111111111111111111111111111111111000000000000000"),
("1111111111111111111111111111111111111111111111111111111100000000000000"),
("1111111111111111111111111111111111111111111111111111111110000000000000"),
("1111111111111111111111111111111111111111111111111111111111000000000000"),
("1111111111111111111111111111111111111111111111111111111111100000000000"),
("1111111111111111111111111111111111111111111111111111111111110000000000"),
("1111111111111111111111111111111111111111111111111111111111111000000000"),
("1111111111111111111111111111111111111111111111111111111111111100000000"),
("1111111111111111111111111111111111111111111111111111111111111110000000"),
("1111111111111111111111111111111111111111111111111111111111111111000000"),
("1111111111111111111111111111111111111111111111111111111111111111100000"),
("1111111111111111111111111111111111111111111111111111111111111111110000"),
("1111111111111111111111111111111111111111111111111111111111111111111000"),
("1111111111111111111111111111111111111111111111111111111111111111111100"),
("1111111111111111111111111111111111111111111111111111111111111111111110"),
("1111111111111111111111111111111111111111111111111111111111111111111111")
);
	
	--left_up_slope:
	constant left_up_slope_start_x 	: integer := 30;
	constant left_up_slope_start_y 	: integer := 30;
	constant left_up_slope_X_size 	: integer := 70;
	constant left_up_slope_Y_size 	: integer := 70;
	constant left_up_slope_color  	: std_logic_vector(7 downto 0) := x"83";
	constant left_up_slope_bounce_type : std_logic_vector(4 downto 0) := left_up_slope;
	signal left_up_slope_end_x : integer;
	signal left_up_slope_end_y : integer;
	signal left_up_slope_drawing_X : std_logic := '0';
	signal left_up_slope_drawing_Y : std_logic := '0';
	signal left_up_slope_drawing_req : std_logic := '0';
	signal left_up_slope_Coord_X : integer := 0;-- offset from start position 
	signal left_up_slope_Coord_Y : integer := 0;
	--/left_up_slope
	
	type left_up_slope_object_form is array (0 to left_up_slope_Y_size - 1 , 0 to left_up_slope_X_size - 1) of std_logic;
	constant left_up_slope_object : left_up_slope_object_form := (
("0111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111110"),
("1111111111111111111111111111111111111111111111111111111111111111111100"),
("1111111111111111111111111111111111111111111111111111111111111111111000"),
("1111111111111111111111111111111111111111111111111111111111111111110000"),
("1111111111111111111111111111111111111111111111111111111111111111100000"),
("1111111111111111111111111111111111111111111111111111111111111111000000"),
("1111111111111111111111111111111111111111111111111111111111111110000000"),
("1111111111111111111111111111111111111111111111111111111111111100000000"),
("1111111111111111111111111111111111111111111111111111111111111000000000"),
("1111111111111111111111111111111111111111111111111111111111110000000000"),
("1111111111111111111111111111111111111111111111111111111111100000000000"),
("1111111111111111111111111111111111111111111111111111111111000000000000"),
("1111111111111111111111111111111111111111111111111111111110000000000000"),
("1111111111111111111111111111111111111111111111111111111100000000000000"),
("1111111111111111111111111111111111111111111111111111111000000000000000"),
("1111111111111111111111111111111111111111111111111111110000000000000000"),
("1111111111111111111111111111111111111111111111111111100000000000000000"),
("1111111111111111111111111111111111111111111111111111000000000000000000"),
("1111111111111111111111111111111111111111111111111110000000000000000000"),
("1111111111111111111111111111111111111111111111111100000000000000000000"),
("1111111111111111111111111111111111111111111111111000000000000000000000"),
("1111111111111111111111111111111111111111111111110000000000000000000000"),
("1111111111111111111111111111111111111111111111100000000000000000000000"),
("1111111111111111111111111111111111111111111111000000000000000000000000"),
("1111111111111111111111111111111111111111111110000000000000000000000000"),
("1111111111111111111111111111111111111111111100000000000000000000000000"),
("1111111111111111111111111111111111111111111000000000000000000000000000"),
("1111111111111111111111111111111111111111110000000000000000000000000000"),
("1111111111111111111111111111111111111111100000000000000000000000000000"),
("1111111111111111111111111111111111111111000000000000000000000000000000"),
("1111111111111111111111111111111111111110000000000000000000000000000000"),
("1111111111111111111111111111111111111100000000000000000000000000000000"),
("1111111111111111111111111111111111111000000000000000000000000000000000"),
("1111111111111111111111111111111111110000000000000000000000000000000000"),
("1111111111111111111111111111111111100000000000000000000000000000000000"),
("1111111111111111111111111111111111000000000000000000000000000000000000"),
("1111111111111111111111111111111110000000000000000000000000000000000000"),
("1111111111111111111111111111111100000000000000000000000000000000000000"),
("1111111111111111111111111111111000000000000000000000000000000000000000"),
("1111111111111111111111111111110000000000000000000000000000000000000000"),
("1111111111111111111111111111100000000000000000000000000000000000000000"),
("1111111111111111111111111111000000000000000000000000000000000000000000"),
("1111111111111111111111111110000000000000000000000000000000000000000000"),
("1111111111111111111111111100000000000000000000000000000000000000000000"),
("1111111111111111111111111000000000000000000000000000000000000000000000"),
("1111111111111111111111110000000000000000000000000000000000000000000000"),
("1111111111111111111111100000000000000000000000000000000000000000000000"),
("1111111111111111111111000000000000000000000000000000000000000000000000"),
("1111111111111111111110000000000000000000000000000000000000000000000000"),
("1111111111111111111100000000000000000000000000000000000000000000000000"),
("1111111111111111111000000000000000000000000000000000000000000000000000"),
("1111111111111111110000000000000000000000000000000000000000000000000000"),
("1111111111111111100000000000000000000000000000000000000000000000000000"),
("1111111111111111000000000000000000000000000000000000000000000000000000"),
("1111111111111110000000000000000000000000000000000000000000000000000000"),
("1111111111111000000000000000000000000000000000000000000000000000000000"),
("1111111111111000000000000000000000000000000000000000000000000000000000"),
("1111111111110000000000000000000000000000000000000000000000000000000000"),
("1111111111100000000000000000000000000000000000000000000000000000000000"),
("1111111110000000000000000000000000000000000000000000000000000000000000"),
("1111111110000000000000000000000000000000000000000000000000000000000000"),
("1111111100000000000000000000000000000000000000000000000000000000000000"),
("1111111000000000000000000000000000000000000000000000000000000000000000"),
("1111100000000000000000000000000000000000000000000000000000000000000000"),
("1111100000000000000000000000000000000000000000000000000000000000000000"),
("1111000000000000000000000000000000000000000000000000000000000000000000"),
("1110000000000000000000000000000000000000000000000000000000000000000000"),
("1100000000000000000000000000000000000000000000000000000000000000000000")
);
	
	--right_down_slope:
	constant right_down_slope_start_x 	: integer := 490;
	constant right_down_slope_start_y 	: integer := 310;
	constant right_down_slope_X_size 	: integer := 70;
	constant right_down_slope_Y_size 	: integer := 70;
	constant right_down_slope_color  	: std_logic_vector(7 downto 0) := x"83";
	constant right_down_slope_bounce_type : std_logic_vector(4 downto 0) := right_down_slope;
	signal right_down_slope_end_x : integer;
	signal right_down_slope_end_y : integer;
	signal right_down_slope_drawing_X : std_logic := '0';
	signal right_down_slope_drawing_Y : std_logic := '0';
	signal right_down_slope_drawing_req : std_logic := '0';
	signal right_down_slope_Coord_X : integer := 0;-- offset from start position 
	signal right_down_slope_Coord_Y : integer := 0;
	--/right_down_slope
	
	type right_down_slope_object_form is array (0 to right_down_slope_Y_size - 1 , 0 to right_down_slope_X_size - 1) of std_logic;
	constant right_down_slope_object : right_down_slope_object_form := (
("0000000000000000000000000000000000000000000000000000000000000000000001"),
("0000000000000000000000000000000000000000000000000000000000000000000011"),
("0000000000000000000000000000000000000000000000000000000000000000000111"),
("0000000000000000000000000000000000000000000000000000000000000000001111"),
("0000000000000000000000000000000000000000000000000000000000000000011111"),
("0000000000000000000000000000000000000000000000000000000000000000111111"),
("0000000000000000000000000000000000000000000000000000000000000001111111"),
("0000000000000000000000000000000000000000000000000000000000000011111111"),
("0000000000000000000000000000000000000000000000000000000000000111111111"),
("0000000000000000000000000000000000000000000000000000000000001111111111"),
("0000000000000000000000000000000000000000000000000000000000011111111111"),
("0000000000000000000000000000000000000000000000000000000000111111111111"),
("0000000000000000000000000000000000000000000000000000000001111111111111"),
("0000000000000000000000000000000000000000000000000000000011111111111111"),
("0000000000000000000000000000000000000000000000000000000111111111111111"),
("0000000000000000000000000000000000000000000000000000001111111111111111"),
("0000000000000000000000000000000000000000000000000000011111111111111111"),
("0000000000000000000000000000000000000000000000000000111111111111111111"),
("0000000000000000000000000000000000000000000000000001111111111111111111"),
("0000000000000000000000000000000000000000000000000011111111111111111111"),
("0000000000000000000000000000000000000000000000000111111111111111111111"),
("0000000000000000000000000000000000000000000000001111111111111111111111"),
("0000000000000000000000000000000000000000000000011111111111111111111111"),
("0000000000000000000000000000000000000000000000111111111111111111111111"),
("0000000000000000000000000000000000000000000001111111111111111111111111"),
("0000000000000000000000000000000000000000000011111111111111111111111111"),
("0000000000000000000000000000000000000000000111111111111111111111111111"),
("0000000000000000000000000000000000000000001111111111111111111111111111"),
("0000000000000000000000000000000000000000011111111111111111111111111111"),
("0000000000000000000000000000000000000000111111111111111111111111111111"),
("0000000000000000000000000000000000000001111111111111111111111111111111"),
("0000000000000000000000000000000000000011111111111111111111111111111111"),
("0000000000000000000000000000000000000111111111111111111111111111111111"),
("0000000000000000000000000000000000001111111111111111111111111111111111"),
("0000000000000000000000000000000000011111111111111111111111111111111111"),
("0000000000000000000000000000000000111111111111111111111111111111111111"),
("0000000000000000000000000000000001111111111111111111111111111111111111"),
("0000000000000000000000000000000011111111111111111111111111111111111111"),
("0000000000000000000000000000000111111111111111111111111111111111111111"),
("0000000000000000000000000000001111111111111111111111111111111111111111"),
("0000000000000000000000000000011111111111111111111111111111111111111111"),
("0000000000000000000000000000111111111111111111111111111111111111111111"),
("0000000000000000000000000001111111111111111111111111111111111111111111"),
("0000000000000000000000000011111111111111111111111111111111111111111111"),
("0000000000000000000000000111111111111111111111111111111111111111111111"),
("0000000000000000000000001111111111111111111111111111111111111111111111"),
("0000000000000000000000011111111111111111111111111111111111111111111111"),
("0000000000000000000000111111111111111111111111111111111111111111111111"),
("0000000000000000000001111111111111111111111111111111111111111111111111"),
("0000000000000000000011111111111111111111111111111111111111111111111111"),
("0000000000000000000111111111111111111111111111111111111111111111111111"),
("0000000000000000001111111111111111111111111111111111111111111111111111"),
("0000000000000000011111111111111111111111111111111111111111111111111111"),
("0000000000000000111111111111111111111111111111111111111111111111111111"),
("0000000000000001111111111111111111111111111111111111111111111111111111"),
("0000000000000011111111111111111111111111111111111111111111111111111111"),
("0000000000000111111111111111111111111111111111111111111111111111111111"),
("0000000000001111111111111111111111111111111111111111111111111111111111"),
("0000000000011111111111111111111111111111111111111111111111111111111111"),
("0000000000111111111111111111111111111111111111111111111111111111111111"),
("0000000001111111111111111111111111111111111111111111111111111111111111"),
("0000000011111111111111111111111111111111111111111111111111111111111111"),
("0000000111111111111111111111111111111111111111111111111111111111111111"),
("0000001111111111111111111111111111111111111111111111111111111111111111"),
("0000011111111111111111111111111111111111111111111111111111111111111111"),
("0000111111111111111111111111111111111111111111111111111111111111111111"),
("0001111111111111111111111111111111111111111111111111111111111111111111"),
("0011111111111111111111111111111111111111111111111111111111111111111111"),
("0111111111111111111111111111111111111111111111111111111111111111111111"),
("1111111111111111111111111111111111111111111111111111111111111111111111")
);

	
	--right_up_slope:
	constant right_up_slope_start_x 	: integer := 540;
--	constant right_up_slope_start_x2 	: integer := 500;
	constant right_up_slope_start_y 	: integer := 30;
	constant right_up_slope_X_size 	: integer := 70;
	constant right_up_slope_Y_size 	: integer := 70;
	constant right_up_slope_color  	: std_logic_vector(7 downto 0) := x"83";
	constant right_up_slope_bounce_type : std_logic_vector(4 downto 0) := right_up_slope;
	signal right_up_slope_end_x : integer;
--	signal right_up_slope_end_x2 : integer;
	signal right_up_slope_end_y : integer;
	signal right_up_slope_drawing_X : std_logic := '0';
--	signal right_up_slope_drawing_X2 : std_logic := '0';
	signal right_up_slope_drawing_Y : std_logic := '0';
	signal right_up_slope_drawing_req : std_logic := '0';
	signal right_up_slope_Coord_X : integer := 0;-- offset from start position 
--	signal right_up_slope_Coord_X2 : integer := 0;-- offset from start position 
	signal right_up_slope_Coord_Y : integer := 0;
	
	constant right_up_slope_begin_offset : integer := -40;
	
	signal right_up_slope_begin_drawing_X : std_logic := '0';
	signal right_up_slope_begin_Coord_X : integer := 0;-- offset from start position 

	--/right_up_slope

	type right_up_slope_object_form is array (0 to right_up_slope_Y_size - 1 , 0 to right_up_slope_X_size - 1) of std_logic;
	constant right_up_slope_object : right_up_slope_object_form := (
("1111111111111111111111111111111111111111111111111111111111111111111111"),
("0111111111111111111111111111111111111111111111111111111111111111111111"),
("0011111111111111111111111111111111111111111111111111111111111111111111"),
("0001111111111111111111111111111111111111111111111111111111111111111111"),
("0000111111111111111111111111111111111111111111111111111111111111111111"),
("0000011111111111111111111111111111111111111111111111111111111111111111"),
("0000001111111111111111111111111111111111111111111111111111111111111111"),
("0000000111111111111111111111111111111111111111111111111111111111111111"),
("0000000011111111111111111111111111111111111111111111111111111111111111"),
("0000000001111111111111111111111111111111111111111111111111111111111111"),
("0000000000111111111111111111111111111111111111111111111111111111111111"),
("0000000000011111111111111111111111111111111111111111111111111111111111"),
("0000000000001111111111111111111111111111111111111111111111111111111111"),
("0000000000000111111111111111111111111111111111111111111111111111111111"),
("0000000000000011111111111111111111111111111111111111111111111111111111"),
("0000000000000001111111111111111111111111111111111111111111111111111111"),
("0000000000000000111111111111111111111111111111111111111111111111111111"),
("0000000000000000011111111111111111111111111111111111111111111111111111"),
("0000000000000000001111111111111111111111111111111111111111111111111111"),
("0000000000000000000111111111111111111111111111111111111111111111111111"),
("0000000000000000000011111111111111111111111111111111111111111111111111"),
("0000000000000000000001111111111111111111111111111111111111111111111111"),
("0000000000000000000000111111111111111111111111111111111111111111111111"),
("0000000000000000000000011111111111111111111111111111111111111111111111"),
("0000000000000000000000001111111111111111111111111111111111111111111111"),
("0000000000000000000000000111111111111111111111111111111111111111111111"),
("0000000000000000000000000011111111111111111111111111111111111111111111"),
("0000000000000000000000000001111111111111111111111111111111111111111111"),
("0000000000000000000000000000111111111111111111111111111111111111111111"),
("0000000000000000000000000000011111111111111111111111111111111111111111"),
("0000000000000000000000000000001111111111111111111111111111111111111111"),
("0000000000000000000000000000000111111111111111111111111111111111111111"),
("0000000000000000000000000000000011111111111111111111111111111111111111"),
("0000000000000000000000000000000001111111111111111111111111111111111111"),
("0000000000000000000000000000000000111111111111111111111111111111111111"),
("0000000000000000000000000000000000011111111111111111111111111111111111"),
("0000000000000000000000000000000000001111111111111111111111111111111111"),
("0000000000000000000000000000000000000111111111111111111111111111111111"),
("0000000000000000000000000000000000000011111111111111111111111111111111"),
("0000000000000000000000000000000000000001111111111111111111111111111111"),
("0000000000000000000000000000000000000000111111111111111111111111111111"),
("0000000000000000000000000000000000000000011111111111111111111111111111"),
("0000000000000000000000000000000000000000001111111111111111111111111111"),
("0000000000000000000000000000000000000000000111111111111111111111111111"),
("0000000000000000000000000000000000000000000011111111111111111111111111"),
("0000000000000000000000000000000000000000000001111111111111111111111111"),
("0000000000000000000000000000000000000000000000111111111111111111111111"),
("0000000000000000000000000000000000000000000000011111111111111111111111"),
("0000000000000000000000000000000000000000000000001111111111111111111111"),
("0000000000000000000000000000000000000000000000000111111111111111111111"),
("0000000000000000000000000000000000000000000000000011111111111111111111"),
("0000000000000000000000000000000000000000000000000001111111111111111111"),
("0000000000000000000000000000000000000000000000000000111111111111111111"),
("0000000000000000000000000000000000000000000000000000011111111111111111"),
("0000000000000000000000000000000000000000000000000000001111111111111111"),
("0000000000000000000000000000000000000000000000000000000111111111111111"),
("0000000000000000000000000000000000000000000000000000000011111111111111"),
("0000000000000000000000000000000000000000000000000000000001111111111111"),
("0000000000000000000000000000000000000000000000000000000000111111111111"),
("0000000000000000000000000000000000000000000000000000000000011111111111"),
("0000000000000000000000000000000000000000000000000000000000001111111111"),
("0000000000000000000000000000000000000000000000000000000000000111111111"),
("0000000000000000000000000000000000000000000000000000000000000011111111"),
("0000000000000000000000000000000000000000000000000000000000000001111111"),
("0000000000000000000000000000000000000000000000000000000000000000111111"),
("0000000000000000000000000000000000000000000000000000000000000000011111"),
("0000000000000000000000000000000000000000000000000000000000000000001111"),
("0000000000000000000000000000000000000000000000000000000000000000000111"),
("0000000000000000000000000000000000000000000000000000000000000000000011"),
("0000000000000000000000000000000000000000000000000000000000000000000001")
);	
	
	
--tunnel_wall:
	constant tunnel_wall_start_x 	: integer := 560;
	constant tunnel_wall_start_y 	: integer := 100;
	constant tunnel_wall_X_size 	: integer := 50;
	constant tunnel_wall_Y_size 	: integer := 350;
	constant tunnel_wall_color  	: std_logic_vector(7 downto 0) := x"d0";
	constant tunnel_wall_bounce_type : std_logic_vector(4 downto 0) := right_vertical_wall;
	signal tunnel_wall_end_x : integer;
	signal tunnel_wall_end_y : integer;
	signal tunnel_wall_drawing_X : std_logic := '0';
	signal tunnel_wall_drawing_Y : std_logic := '0';
	signal tunnel_wall_drawing_req : std_logic := '0';
	signal tunnel_wall_Coord_X : integer := 0;-- offset from start position 
	signal tunnel_wall_Coord_Y : integer := 0;
--/tunnel_wall
	
	type tunnel_wall_object_form is array (0 to tunnel_wall_Y_size - 1 , 0 to tunnel_wall_X_size - 1) of std_logic;
	constant tunnel_wall_object : tunnel_wall_object_form := (
("00000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111110000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111"),
("11111111111111111111111111111111111111111111111111")
);	



--stage_left:
	constant stage_left_start_x 	: integer := 30;
	constant stage_left_start_y 	: integer := 380;
	constant stage_left_X_size 	: integer := 190;
	constant stage_left_Y_size 	: integer := 70;
	constant stage_left_color  	: std_logic_vector(7 downto 0) := x"d0";
	constant stage_left_bounce_type1 : std_logic_vector(4 downto 0) := horizontal_floor;
	constant stage_left_bounce_type2 : std_logic_vector(4 downto 0) := left_vertical_wall;
	signal stage_left_end_x : integer;
	signal stage_left_end_y : integer;
	signal stage_left_drawing_X : std_logic := '0';
	signal stage_left_drawing_Y : std_logic := '0';
	signal stage_left_drawing_req : std_logic := '0';
--/stage_left

 --stage_right:
	constant stage_right_start_x 	: integer := 380;
	constant stage_right_start_y 	: integer := 380;
	constant stage_right_X_size 	: integer := 180;
	constant stage_right_Y_size 	: integer := 70;
	constant stage_right_color  	: std_logic_vector(7 downto 0) := x"d0";
	constant stage_right_bounce_type1 : std_logic_vector(4 downto 0) := horizontal_floor;
	constant stage_right_bounce_type2 : std_logic_vector(4 downto 0) := right_vertical_wall;
	signal stage_right_end_x : integer;
	signal stage_right_end_y : integer;
	signal stage_right_drawing_X : std_logic := '0';
	signal stage_right_drawing_Y : std_logic := '0';
	signal stage_right_drawing_req : std_logic := '0';
--/stage_right


 --start_message:
	constant start_message_start_x 	: integer := 200;
	constant start_message_start_y 	: integer := 280;
	constant start_message_X_size 	: integer := 200;
	constant start_message_Y_size 	: integer := 100;
	constant start_message_color  	: std_logic_vector(7 downto 0) := x"ff";
	constant start_message_bounce_type : std_logic_vector(4 downto 0) := no_bounce;
	signal start_message_end_x : integer;
	signal start_message_end_y : integer;
	signal start_message_drawing_X : std_logic := '0';
	signal start_message_drawing_Y : std_logic := '0';
	signal start_message_drawing_req : std_logic := '0';
	signal start_message_Coord_X : integer := 0;-- offset from start position 
	signal start_message_Coord_Y : integer := 0;
--/start_message

type start_message_object_form is array (0 to start_message_Y_size - 1 , 0 to start_message_X_size - 1) of std_logic;
constant start_message_object : start_message_object_form := (
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00001111111111000001111111111000000111111111111000001111111000000001111111000000000000000111111000000111111111000000000111000000000000111111000000011111111111100000011111111111111000000111111000000000"),
("00001111111111100001111111111110000111111111111100011111111100000011111111100000000000001111111110000111111111110000000111100000000001111111110000011111111111100000011111111111111100001111111110000000"),
("00001111111111110001111111111111000111111111111100111111111110000111111111110000000000011111111110000111111111111000000111100000000011111111111000011111111111100000011111111111111100011111111111000000"),
("00001111111111111001111111111111000111111111111000111111111110000111111111110000000000111111111111000111111111111100001111100000000111111111111000011111111111100000011111111111111000111111111111000000"),
("00001110000001111001111000000111100111000000000001111000001111001111000001111000000000111100001111000111000001111100001111110000000111100001111100011100000000000000000000011100000001111100001111100000"),
("00001110000000111001111000000111100111000000000001111000001111001111000001111000000000111000000111000111000000011100001111110000001111000000111100011100000000000000000000011100000001111000000111100000"),
("00001110000000111101111000000011100111000000000001110000000111001110000000111000000000111000000111100111000000011100001111110000001110000000011100011100000000000000000000011100000001110000000011110000"),
("00001110000000111101111000000011100111000000000001110000000111001110000000111000000000111000000111100111000000011100011101110000001110000000011110011100000000000000000000011100000011110000000011110000"),
("00001110000000111101111000000011100111000000000001110000000111001110000000111000000000111000000011100111000000011100011101111000011110000000011100011100000000000000000000011100000011110000000001110000"),
("00001110000000111101111000000011100111000000000001111000000000001111000000000000000000111000000000000111000000011100011100111000011110000000000000011100000000000000000000011100000011100000000001110000"),
("00001110000000111101111000000011100111000000000001111100000000001111100000000000000000111110000000000111000000011100011100111000011100000000000000011100000000000000000000011100000011100000000001110000"),
("00001110000000111001110000000111100111111111110000111111100000000111111100000000000000111111100000000111000000111100111100111000011100000000000000011111111111000000000000011100000011100000000001111000"),
("00001111000001111001111111111111000111111111111000111111111000000111111111000000000000011111111100000111000001111100111000111100011100000000000000011111111111000000000000011100000011100000000001111000"),
("00001111111111111001111111111111000111111111111000011111111110000011111111110000000000001111111110000111111111111100111000111100011100000000000000011111111111000000000000011100000011100000000001111000"),
("00001111111111110001111111111110000111111111111000000111111110000000111111111000000000000111111111000111111111111000111000011100011100000000000000011111111111000000000000011100000011100000000001111000"),
("00001111111111100001111111111111000111000000000000000001111111000000001111111000000000000000111111100111111111110001111000011100011100000000000000011100000000000000000000011100000011100000000001111000"),
("00001111111111000001111000001111000111000000000000000000001111000000000001111100000000000000001111100111111111100001111111111110011100000000001100011100000000000000000000011100000011100000000001111000"),
("00001110000000000001111000000111100111000000000000000000000111100000000000111100000000000000000111100111000000000001111111111110011100000000011110011100000000000000000000011100000011100000000001110000"),
("00001110000000000001111000000111100111000000000011110000000111101110000000111100000001110000000011100111000000000001111111111110011110000000011110011100000000000000000000011100000011100000000001110000"),
("00001110000000000001111000000011100111000000000011110000000011101110000000011100000001110000000011100111000000000011111111111110011110000000011110011100000000000000000000011100000011110000000001110000"),
("00001110000000000001111000000011100111000000000001110000000011101110000000011100000001110000000011100111000000000011100000001111001110000000011100011100000000000000000000011100000011110000000011110000"),
("00001110000000000001111000000011100111000000000001110000000111101110000000111100000001111000000011100111000000000011100000001111001111000000011100011100000000000000000000011100000001111000000011100000"),
("00001110000000000001111000000011100111000000000001111000000111101111000000111100000001111000000111100111000000000011100000000111001111000000111100011100000000000000000000011100000001111000000111100000"),
("00001110000000000001111000000011100111111111111001111100001111001111100001111000000000111100001111100111000000000111100000000111000111100001111000011111111111100000000000011100000000111100001111100000"),
("00001110000000000001111000000011100111111111111100111111111111000111111111111000000000111111111111000111000000000111100000000111100111111111111000011111111111100000000000011100000000111111111111000000"),
("00001110000000000001111000000011100111111111111100111111111110000011111111110000000000011111111111000111000000000111000000000111100011111111110000011111111111100000000000011100000000011111111110000000"),
("00001110000000000001111000000011110111111111111100001111111100000001111111100000000000001111111110000111000000000111000000000111100001111111100000011111111111100000000000011100000000001111111100000000"),
("00000000000000000000000000000000000000000000000000000111110000000000111110000000000000000011111000000000000000000000000000000000000000011111000000000000000000000000000000000000000000000011111000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000011111100000111111111111100000110000000011111111000000111111111111100000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000111111110001111111111111100001110000000111111111111001111111111111100000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000001111111111001111111111111100011111000000111111111111101111111111111100000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000011111111111001111111111111100011111000000111111111111101111111111111100000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000011110000111100111011110111100011111000000111100001111110101011110111000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000111100000011100000001110000000011111000000111100000011110000001110000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000111100000011100000001110000000111111100000111100000001110000001110000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000111100000011100000001110000000111011100000111100000001110000001110000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000111100000011100000001110000000111011100000111100000001110000001110000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000111100000000000000001110000000111011100000111100000001110000001110000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000111110000000000000001110000001111011110000111100000001110000001110000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000011111100000000000001110000001110001110000111100000011110000001110000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000011111111100000000001110000001110001110000111100001111100000001110000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000001111111111000000001110000001110001110000111111111111100000001110000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000011111111100000001110000011110001111000111111111111000000001110000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000111111100000001110000011100000111000111111111111100000001110000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000111110000001110000011111111111000111100000111100000001110000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000011110000001110000011111111111000111100000011110000001110000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000111000000001110000001110000111111111111100111100000011110000001110000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000111000000001110000001110000111111111111100111100000001110000001110000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000111000000001110000001110000111000000011100111100000001110000001110000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000111000000001110000001110000111000000011100111100000001110000001110000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000111100000011110000001110001111000000011110111100000001110000001110000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000011110000011110000001110001110000000011110111100000001110000001110000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000011111111111100000001110001110000000001110111100000001110000001110000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000001111111111100000001110001110000000001110111100000001110000001110000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000111111111000000001110011110000000001111111100000001111000001110000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000011111100000000001100001100000000000110011000000000110000001100000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000")
);





------------------------------- obsticle -------------------------------------------------------------------

 --game_over_message:
	constant game_over_message_start_x 	: integer := 200;
	constant game_over_message_start_y 	: integer := 280;
	constant game_over_message_X_size 	: integer := 200;
	constant game_over_message_Y_size 	: integer := 100;
	constant game_over_message_color  	: std_logic_vector(7 downto 0) := x"ff";
	constant game_over_message_bounce_type : std_logic_vector(4 downto 0) := no_bounce;
	signal game_over_message_end_x : integer;
	signal game_over_message_end_y : integer;
	signal game_over_message_drawing_X : std_logic := '0';
	signal game_over_message_drawing_Y : std_logic := '0';
	signal game_over_message_drawing_req : std_logic := '0';
	signal game_over_message_Coord_X : integer := 0;-- offset from start position 
	signal game_over_message_Coord_Y : integer := 0;
--/game_over_message

type game_over_message_object_form is array (0 to game_over_message_Y_size - 1 , 0 to game_over_message_X_size - 1) of std_logic;
constant game_over_message_object : game_over_message_object_form := (
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000111111111100000000000000011111000000000011111000000000000001111100001111111111111111100000000000000000111111111100000001111000000000000111110111111111111111110001111111111111100000000000"),
("00000000000001111111111111000000000000011111000000000011111000000000000011111100001111111111111111100000000000000011111111111110000001111100000000000111110111111111111111110001111111111111111000000000"),
("00000000000111111111111111100000000000111111000000000011111100000000000011111100001111111111111111100000000000000111111111111111000001111100000000000111100111111111111111110001111111111111111100000000"),
("00000000000111111111111111100000000000111111100000000011111100000000000011111100001111111111111111100000000000001111111111111111100000111100000000000111100111111111111111110001111111111111111110000000"),
("00000000001111110000001111110000000000111111100000000011111100000000000111111100001111000000000000000000000000001111110000001111110000111100000000001111100111100000000000000001111000000001111110000000"),
("00000000011111100000000011111000000001111111100000000011111110000000000111111100001111000000000000000000000000011111000000000111110000111110000000001111000111100000000000000001111000000000011110000000"),
("00000000011111000000000011111000000001111011110000000011111110000000000111111100001111000000000000000000000000011111000000000011111000111110000000001111000111100000000000000001111000000000011111000000"),
("00000000011110000000000001111000000001111011110000000011111110000000001111111100001111000000000000000000000000111110000000000001111000011110000000011111000111100000000000000001111000000000011111000000"),
("00000000111110000000000001111000000001111011110000000011111111000000001111111100001111000000000000000000000000111100000000000001111100011110000000011111000111100000000000000001111000000000011111000000"),
("00000000111100000000000001111000000011110011111000000011111111000000001111111100001111000000000000000000000000111100000000000001111100011111000000011110000111100000000000000001111000000000011111000000"),
("00000000111100000000000000000000000011110001111000000011111111000000011110111100001111000000000000000000000000111100000000000000111100001111000000011110000111100000000000000001111000000000011110000000"),
("00000000111100000000000000000000000011110001111000000011110111100000011110111100001111000000000000000000000001111100000000000000111100001111000000111110000111100000000000000001111000000000011110000000"),
("00000001111100000000000000000000000111100001111100000011110111100000011110111100001111111111111111000000000001111100000000000000111100001111100000111100000111111111111111100001111000000001111110000000"),
("00000001111100000001111111111000000111100000111100000011110111100000011110111100001111111111111111000000000001111000000000000000111100001111100000111100000111111111111111100001111111111111111100000000"),
("00000001111100000011111111111100000111100000111100000011110011110000111100111100001111111111111111000000000001111000000000000000111100000111100000111100000111111111111111100001111111111111111000000000"),
("00000001111100000011111111111100001111000000111110000011110011110000111100111100001111111111111111000000000001111000000000000000111100000111100001111000000111111111111111100001111111111111111000000000"),
("00000001111100000011111111111100001111111111111110000011110011110000111100111100001111000000000000000000000001111000000000000000111100000111110001111000000111100000000000000001111111111111111100000000"),
("00000001111100000001111111111100001111111111111110000011110001110001111000111100001111000000000000000000000001111100000000000000111100000011110001111000000111100000000000000001111000000001111100000000"),
("00000000111100000000000000111100011111111111111111000011110001111001111000111100001111000000000000000000000001111100000000000000111100000011110011111000000111100000000000000001111000000000111110000000"),
("00000000111100000000000000111100011111111111111111000011110001111001111000111100001111000000000000000000000000111100000000000000111100000011110011110000000111100000000000000001111000000000011110000000"),
("00000000111110000000000001111100011111111111111111000011110001111011110000111100001111000000000000000000000000111100000000000001111100000001111011110000000111100000000000000001111000000000011110000000"),
("00000000111110000000000001111100111110000000001111100011110000111111110000111100001111000000000000000000000000111110000000000001111000000001111011110000000111100000000000000001111000000000011110000000"),
("00000000011111000000000011111100111100000000001111100011110000111111110000111100001111000000000000000000000000011110000000000011111000000001111111100000000111100000000000000001111000000000011110000000"),
("00000000011111000000000011111100111100000000000111100011110000111111100000111100001111000000000000000000000000011111000000000111111000000001111111100000000111100000000000000001111000000000011110000000"),
("00000000001111100000001111111101111100000000000111100011110000011111100000111100001111000000000000000000000000001111100000001111110000000000111111100000000111100000000000000001111000000000011110000000"),
("00000000001111111100111111111101111000000000000111110011110000011111100000111100001111111111111111100000000000001111111100111111100000000000111111100000000111111111111111110001111000000000011110000000"),
("00000000000111111111111111111101111000000000000111110011110000011111100000111100001111111111111111100000000000000111111111111111000000000000111111000000000111111111111111110001111000000000011111000000"),
("00000000000011111111111110111111111000000000000011110011110000001111000000111100001111111111111111100000000000000011111111111110000000000000011111000000000111111111111111110001111000000000011111000000"),
("00000000000000111111111100011011111000000000000011111011110000001111000000111100001111111111111111100000000000000000111111111100000000000000011111000000000111111111111111110001111000000000001111000000"),
("00000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000011111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000011110000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000")
);



-- obsticle_up
	constant obsticle_up_start_x 	: integer := 150;
	constant obsticle_up_start_y 	: integer := 100;
	constant obsticle_up_X_size 	: integer := 20;
	constant obsticle_up_Y_size 	: integer := 20;
	constant obsticle_up_color  	: std_logic_vector(7 downto 0) := x"e1";
	constant obsticle_up_bounce_type : std_logic_vector(4 downto 0) := horizontal_floor;
	signal obsticle_up_end_x : integer;
	signal obsticle_up_end_y : integer;
	signal obsticle_up_drawing_X : std_logic := '0';
	signal obsticle_up_drawing_Y : std_logic := '0';
	signal obsticle_up_drawing_req : std_logic := '0';
--/obsticle_up


-- obsticle_left_up
	constant obsticle_left_up_start_x 	: integer := 130;
	constant obsticle_left_up_start_y 	: integer := 100;
	constant obsticle_left_up_X_size 	: integer := 20;
	constant obsticle_left_up_Y_size 	: integer := 20;
	constant obsticle_left_up_color  	: std_logic_vector(7 downto 0) := x"ff";
	constant obsticle_left_up_bounce_type : std_logic_vector(4 downto 0) := right_down_slope;
	signal obsticle_left_up_end_x : integer;
	signal obsticle_left_up_end_y : integer;
	signal obsticle_left_up_drawing_X : std_logic := '0';
	signal obsticle_left_up_drawing_Y : std_logic := '0';
	signal obsticle_left_up_drawing_req : std_logic := '0';
	signal obsticle_left_up_Coord_X : integer := 0;-- offset from start position 
	signal obsticle_left_up_Coord_Y : integer := 0;

--/obsticle_left_up

-- obsticle_left
	constant obsticle_left_start_x 	: integer := 130;
	constant obsticle_left_start_y 	: integer := 120;
	constant obsticle_left_X_size 	: integer := 30;
	constant obsticle_left_Y_size 	: integer := 20;
	constant obsticle_left_color  	: std_logic_vector(7 downto 0) := x"e1";
	constant obsticle_left_bounce_type : std_logic_vector(4 downto 0) := left_vertical_wall;
	signal obsticle_left_end_x : integer;
	signal obsticle_left_end_y : integer;
	signal obsticle_left_drawing_X : std_logic := '0';
	signal obsticle_left_drawing_Y : std_logic := '0';
	signal obsticle_left_drawing_req : std_logic := '0';
--/obsticle_left


-- obsticle_left_down
	constant obsticle_left_down_start_x 	: integer := 130;
	constant obsticle_left_down_start_y 	: integer := 140;
	constant obsticle_left_down_X_size 	: integer := 20;
	constant obsticle_left_down_Y_size 	: integer := 20;
	constant obsticle_left_down_color  	: std_logic_vector(7 downto 0) := x"ff";
	constant obsticle_left_down_bounce_type : std_logic_vector(4 downto 0) := right_up_slope;
	signal obsticle_left_down_end_x : integer;
	signal obsticle_left_down_end_y : integer;
	signal obsticle_left_down_drawing_X : std_logic := '0';
	signal obsticle_left_down_drawing_Y : std_logic := '0';
	signal obsticle_left_down_drawing_req : std_logic := '0';
	signal obsticle_left_down_Coord_X : integer := 0;-- offset from start position 
	signal obsticle_left_down_Coord_Y : integer := 0;


--/obsticle_left_down

-- obsticle_down
	constant obsticle_down_start_x 	: integer := 150;
	constant obsticle_down_start_y 	: integer := 140;
	constant obsticle_down_X_size 	: integer := 20;
	constant obsticle_down_Y_size 	: integer := 20;
	constant obsticle_down_color  	: std_logic_vector(7 downto 0) := x"e1";
	constant obsticle_down_bounce_type : std_logic_vector(4 downto 0) := horizontal_ceiling;
	signal obsticle_down_end_x : integer;
	signal obsticle_down_end_y : integer;
	signal obsticle_down_drawing_X : std_logic := '0';
	signal obsticle_down_drawing_Y : std_logic := '0';
	signal obsticle_down_drawing_req : std_logic := '0';
--/obsticle_down

-- obsticle_right_down
	constant obsticle_right_down_start_x 	: integer := 170;
	constant obsticle_right_down_start_y 	: integer := 140;
	constant obsticle_right_down_X_size 	: integer := 20;
	constant obsticle_right_down_Y_size 	: integer := 20;
	constant obsticle_right_down_color  	: std_logic_vector(7 downto 0) := x"ff";
	constant obsticle_right_down_bounce_type : std_logic_vector(4 downto 0) := left_up_slope;
	signal obsticle_right_down_end_x : integer;
	signal obsticle_right_down_end_y : integer;
	signal obsticle_right_down_drawing_X : std_logic := '0';
	signal obsticle_right_down_drawing_Y : std_logic := '0';
	signal obsticle_right_down_drawing_req : std_logic := '0';
	signal obsticle_right_down_Coord_X : integer := 0;-- offset from start position 
	signal obsticle_right_down_Coord_Y : integer := 0;


--/obsticle_right_down



-- obsticle_right
	constant obsticle_right_start_x 	: integer := 160;
	constant obsticle_right_start_y 	: integer := 120;
	constant obsticle_right_X_size 	: integer := 30;
	constant obsticle_right_Y_size 	: integer := 20;
	constant obsticle_right_color  	: std_logic_vector(7 downto 0) := x"e1";
	constant obsticle_right_bounce_type : std_logic_vector(4 downto 0) := right_vertical_wall;
	signal obsticle_right_end_x : integer;
	signal obsticle_right_end_y : integer;
	signal obsticle_right_drawing_X : std_logic := '0';
	signal obsticle_right_drawing_Y : std_logic := '0';
	signal obsticle_right_drawing_req : std_logic := '0';
--/obsticle_right



-- obsticle_right_up

	constant obsticle_right_up_start_x 	: integer := 170;
	constant obsticle_right_up_start_y 	: integer := 100;
	constant obsticle_right_up_X_size 	: integer := 20;
	constant obsticle_right_up_Y_size 	: integer := 20;
	constant obsticle_right_up_color  	: std_logic_vector(7 downto 0) := x"ff";
	constant obsticle_right_up_bounce_type : std_logic_vector(4 downto 0) := left_down_slope;
	signal obsticle_right_up_end_x : integer;
	signal obsticle_right_up_end_y : integer;
	signal obsticle_right_up_drawing_X : std_logic := '0';
	signal obsticle_right_up_drawing_Y : std_logic := '0';
	signal obsticle_right_up_drawing_req : std_logic := '0';
	signal obsticle_right_up_Coord_X : integer := 0;-- offset from start position 
	signal obsticle_right_up_Coord_Y : integer := 0;

--/obsticle_right_up


type obsticle_array is array (0 to obsticle_left_up_Y_size - 1 , 0 to obsticle_left_up_X_size - 1) of std_logic;


	constant obsticle_left_up_mask : obsticle_array :=  (
		("00000000000000000001"),
		("00000000000000000011"),
		("00000000000000000111"),
		("00000000000000001111"),
		("00000000000000011111"),
		("00000000000000111111"),
		("00000000000001111111"),
		("00000000000011111111"),
		("00000000000111111111"),
		("00000000001111111111"),
		("00000000011111111111"),
		("00000000111111111111"),
		("00000001111111111111"),
		("00000011111111111111"),
		("00000111111111111111"),
		("00001111111111111111"),
		("00011111111111111111"),
		("00111111111111111111"),
		("01111111111111111111"),
		("11111111111111111111")
		);
	
	
	constant obsticle_left_down_mask : obsticle_array := (
		("11111111111111111111"),
		("01111111111111111111"),
		("00111111111111111111"),
		("00011111111111111111"),
		("00001111111111111111"),
		("00000111111111111111"),
		("00000011111111111111"),
		("00000001111111111111"),
		("00000000111111111111"),
		("00000000011111111111"),
		("00000000001111111111"),
		("00000000000111111111"),
		("00000000000011111111"),
		("00000000000001111111"),
		("00000000000000111111"),
		("00000000000000011111"),
		("00000000000000001111"),
		("00000000000000000111"),
		("00000000000000000011"),
		("00000000000000000001")
		);
	
		
	constant obsticle_right_down_mask : obsticle_array :=  (
		("11111111111111111111"),
		("11111111111111111110"),
		("11111111111111111100"),
		("11111111111111111000"),
		("11111111111111110000"),
		("11111111111111100000"),
		("11111111111111000000"),
		("11111111111110000000"),
		("11111111111100000000"),
		("11111111111000000000"),
		("11111111110000000000"),
		("11111111100000000000"),
		("11111111000000000000"),
		("11111110000000000000"),
		("11111100000000000000"),
		("11111000000000000000"),
		("11110000000000000000"),
		("11100000000000000000"),
		("11000000000000000000"),
		("10000000000000000000")
		);


	constant obsticle_right_up_mask : obsticle_array :=  (
		("10000000000000000000"),
		("11000000000000000000"),
		("11100000000000000000"),
		("11110000000000000000"),
		("11111000000000000000"),
		("11111100000000000000"),
		("11111110000000000000"),
		("11111111000000000000"),
		("11111111100000000000"),
		("11111111110000000000"),
		("11111111111000000000"),
		("11111111111100000000"),
		("11111111111110000000"),
		("11111111111111000000"),
		("11111111111111100000"),
		("11111111111111110000"),
		("11111111111111111000"),
		("11111111111111111100"),
		("11111111111111111110"),
		("11111111111111111111")
		);
	
	constant obsticle_2_x_offset : integer := 100;
	constant obsticle_2_y_offset : integer := 50;
	
-- obsticle_up
	signal obsticle_2_up_drawing_X : std_logic := '0';
	signal obsticle_2_up_drawing_Y : std_logic := '0';
	
--/obsticle_up


-- obsticle_left_up
	signal obsticle_2_left_up_drawing_X : std_logic := '0';
	signal obsticle_2_left_up_drawing_Y : std_logic := '0';
	signal obsticle_2_left_up_Coord_X : integer := 0;-- offset from start position 
	signal obsticle_2_left_up_Coord_Y : integer := 0;

--/obsticle_left_up

-- obsticle_left
	signal obsticle_2_left_drawing_X : std_logic := '0';
	signal obsticle_2_left_drawing_Y : std_logic := '0';
	
--/obsticle_left


-- obsticle_left_down
	signal obsticle_2_left_down_drawing_X : std_logic := '0';
	signal obsticle_2_left_down_drawing_Y : std_logic := '0';
	signal obsticle_2_left_down_Coord_X : integer := 0;-- offset from start position 
	signal obsticle_2_left_down_Coord_Y : integer := 0;


--/obsticle_left_down

-- obsticle_down
	signal obsticle_2_down_drawing_X : std_logic := '0';
	signal obsticle_2_down_drawing_Y : std_logic := '0';
	
--/obsticle_down

-- obsticle_right_down
	signal obsticle_2_right_down_drawing_X : std_logic := '0';
	signal obsticle_2_right_down_drawing_Y : std_logic := '0';
	signal obsticle_2_right_down_Coord_X : integer := 0;-- offset from start position 
	signal obsticle_2_right_down_Coord_Y : integer := 0;


--/obsticle_right_down



-- obsticle_right
	signal obsticle_2_right_drawing_X : std_logic := '0';
	signal obsticle_2_right_drawing_Y : std_logic := '0';
--/obsticle_right



-- obsticle_right_up

	signal obsticle_2_right_up_drawing_X : std_logic := '0';
	signal obsticle_2_right_up_drawing_Y : std_logic := '0';
	signal obsticle_2_right_up_Coord_X : integer := 0;-- offset from start position 
	signal obsticle_2_right_up_Coord_Y : integer := 0;

--/obsticle_right_up


	constant obsticle_3_x_offset : integer := 240;
	constant obsticle_3_y_offset : integer := 50;
	
-- obsticle_up
	signal obsticle_3_up_drawing_X : std_logic := '0';
	signal obsticle_3_up_drawing_Y : std_logic := '0';
	
--/obsticle_up


-- obsticle_left_up
	signal obsticle_3_left_up_drawing_X : std_logic := '0';
	signal obsticle_3_left_up_drawing_Y : std_logic := '0';
	signal obsticle_3_left_up_Coord_X : integer := 0;-- offset from start position 
	signal obsticle_3_left_up_Coord_Y : integer := 0;

--/obsticle_left_up

-- obsticle_left
	signal obsticle_3_left_drawing_X : std_logic := '0';
	signal obsticle_3_left_drawing_Y : std_logic := '0';
	
--/obsticle_left


-- obsticle_left_down
	signal obsticle_3_left_down_drawing_X : std_logic := '0';
	signal obsticle_3_left_down_drawing_Y : std_logic := '0';
	signal obsticle_3_left_down_Coord_X : integer := 0;-- offset from start position 
	signal obsticle_3_left_down_Coord_Y : integer := 0;


--/obsticle_left_down

-- obsticle_down
	signal obsticle_3_down_drawing_X : std_logic := '0';
	signal obsticle_3_down_drawing_Y : std_logic := '0';
	
--/obsticle_down

-- obsticle_right_down
	signal obsticle_3_right_down_drawing_X : std_logic := '0';
	signal obsticle_3_right_down_drawing_Y : std_logic := '0';
	signal obsticle_3_right_down_Coord_X : integer := 0;-- offset from start position 
	signal obsticle_3_right_down_Coord_Y : integer := 0;


--/obsticle_right_down



-- obsticle_right
	signal obsticle_3_right_drawing_X : std_logic := '0';
	signal obsticle_3_right_drawing_Y : std_logic := '0';
--/obsticle_right



-- obsticle_right_up

	signal obsticle_3_right_up_drawing_X : std_logic := '0';
	signal obsticle_3_right_up_drawing_Y : std_logic := '0';
	signal obsticle_3_right_up_Coord_X : integer := 0;-- offset from start position 
	signal obsticle_3_right_up_Coord_Y : integer := 0;

--/obsticle_right_up
------------------------------- /obsticle -------------------------------------------------------------------


	

--		


begin

	-- Calculate objects end boundaries
	left_down_slope_end_x	<= left_down_slope_X_size + left_down_slope_start_x;
	left_down_slope_end_y	<= left_down_slope_Y_size + left_down_slope_start_y;
	
	left_up_slope_end_x	<= left_up_slope_X_size + left_up_slope_start_x;
	left_up_slope_end_y	<= left_up_slope_Y_size + left_up_slope_start_y;
	
	right_down_slope_end_x	<= right_down_slope_X_size + right_down_slope_start_x;
	right_down_slope_end_y	<= right_down_slope_Y_size + right_down_slope_start_y;
	
	right_up_slope_end_x	<= right_up_slope_X_size + right_up_slope_start_x;
	right_up_slope_end_y	<= right_up_slope_Y_size + right_up_slope_start_y;
	
	--right_up_slope_end_x2<= right_up_slope_X_size + right_up_slope_start_x2;
	
	tunnel_wall_end_x	<= tunnel_wall_X_size + tunnel_wall_start_x;
	tunnel_wall_end_y	<= tunnel_wall_Y_size + tunnel_wall_start_y;
	
	stage_left_end_x	<= stage_left_X_size + stage_left_start_x;
	stage_left_end_y	<= stage_left_Y_size + stage_left_start_y;
	
	stage_right_end_x	<= stage_right_X_size + stage_right_start_x;
	stage_right_end_y	<= stage_right_Y_size + stage_right_start_y;
	
	start_message_end_x	<= start_message_X_size + start_message_start_x;
	start_message_end_y	<= start_message_Y_size + start_message_start_y;
	
	game_over_message_end_x	<= game_over_message_X_size + game_over_message_start_x;
	game_over_message_end_y	<= game_over_message_Y_size + game_over_message_start_y;
	
	
	---------------------------------------------------------------
	
	
	floor_end_x	<= floor_X_size + floor_start_x;
	floor_end_y	<= floor_Y_size + floor_start_y;
	
	ceiling_end_x	<= ceiling_X_size + ceiling_start_x;
	ceiling_end_y	<= ceiling_Y_size + ceiling_start_y;
	
	left_wall_end_x	<= left_wall_X_size + left_wall_start_x;
	left_wall_end_y	<= left_wall_Y_size + left_wall_start_y;
	
	right_wall_end_x	<= right_wall_X_size + right_wall_start_x;
	right_wall_end_y	<= right_wall_Y_size + right_wall_start_y;
	
	------ Signals if the game started or if we fell to the pit  -------------------------------------------
	--game_started <= '1' when (oCoord_X  <  game_started_X_bound) else '0';
	--fell_to_pit <= '1' when  (oCoord_X > fell_to_pit_right_X_bound ) and  (oCoord_X < fell_to_pit_right_X_bound ) and  (oCoord_Y > fell_to_pit_upper_Y_bound) else '0';
	
	------------------------------------------------------------------
	
	obsticle_up_end_x <= obsticle_up_X_size + obsticle_up_start_x;
	obsticle_up_end_y <= obsticle_up_Y_size + obsticle_up_start_Y;
	
	obsticle_left_up_end_x <= obsticle_left_up_X_size + obsticle_left_up_start_x;
	obsticle_left_up_end_y <= obsticle_left_up_Y_size + obsticle_left_up_start_Y;
	
	obsticle_left_end_x <= obsticle_left_X_size + obsticle_left_start_x;
	obsticle_left_end_y <= obsticle_left_Y_size + obsticle_left_start_Y;

	obsticle_left_down_end_x <= obsticle_left_down_X_size + obsticle_left_down_start_x;
	obsticle_left_down_end_y <= obsticle_left_down_Y_size + obsticle_left_down_start_Y;

	obsticle_down_end_x <= obsticle_down_X_size + obsticle_down_start_x;
	obsticle_down_end_y <= obsticle_down_Y_size + obsticle_down_start_Y;

	obsticle_right_down_end_x <= obsticle_right_down_X_size + obsticle_right_down_start_x;
	obsticle_right_down_end_y <= obsticle_right_down_Y_size + obsticle_right_down_start_Y;

	obsticle_right_end_x <= obsticle_right_X_size + obsticle_right_start_x;
	obsticle_right_end_y <= obsticle_right_Y_size + obsticle_right_start_Y;

	obsticle_right_up_end_x <= obsticle_right_up_X_size + obsticle_right_up_start_x;
	obsticle_right_up_end_y <= obsticle_right_up_Y_size + obsticle_right_up_start_Y;


	----------------------------------------------------------------------------------
	
	-- test if ooCoord is in the rectangle defined by Start and End 
   floor_drawing_X	<= '1' when  (oCoord_X  >= floor_start_x) and  (oCoord_X < floor_end_x) else '0';
   floor_drawing_Y	<= '1' when  (oCoord_Y  >= floor_start_y) and  (oCoord_Y < floor_end_y) else '0';
	
   ceiling_drawing_X	<= '1' when  (oCoord_X  >= ceiling_start_x) and  (oCoord_X < ceiling_end_x) else '0';
   ceiling_drawing_Y	<= '1' when  (oCoord_Y  >= ceiling_start_y) and  (oCoord_Y < ceiling_end_y) else '0';
	
   left_wall_drawing_X	<= '1' when  (oCoord_X  >= left_wall_start_x) and  (oCoord_X < left_wall_end_x) else '0';
   left_wall_drawing_Y	<= '1' when  (oCoord_Y  >= left_wall_start_y) and  (oCoord_Y < left_wall_end_y) else '0';
	
   right_wall_drawing_X	<= '1' when  (oCoord_X  >= right_wall_start_x) and  (oCoord_X < right_wall_end_x) else '0';
   right_wall_drawing_Y	<= '1' when  (oCoord_Y  >= right_wall_start_y) and  (oCoord_Y < right_wall_end_y) else '0';	
	--------------------------------------------------------------------------------------------------------
	
   left_down_slope_drawing_X	<= '1' when  (oCoord_X  >= left_down_slope_start_x) and  (oCoord_X < left_down_slope_end_x) else '0';
   left_down_slope_drawing_Y	<= '1' when  (oCoord_Y  >= left_down_slope_start_y) and  (oCoord_Y < left_down_slope_end_y) else '0';
	
   left_up_slope_drawing_X	<= '1' when  (oCoord_X  >= left_up_slope_start_x) and  (oCoord_X < left_up_slope_end_x) else '0';
   left_up_slope_drawing_Y	<= '1' when  (oCoord_Y  >= left_up_slope_start_y) and  (oCoord_Y < left_up_slope_end_y) else '0';
	
   right_down_slope_drawing_X	<= '1' when  (oCoord_X  >= right_down_slope_start_x) and  (oCoord_X < right_down_slope_end_x) else '0';
   right_down_slope_drawing_Y	<= '1' when  (oCoord_Y  >= right_down_slope_start_y) and  (oCoord_Y < right_down_slope_end_y) else '0';
	
   right_up_slope_drawing_X	<= '1' when  (oCoord_X  >= right_up_slope_start_x) and  (oCoord_X < right_up_slope_end_x) else '0';
   right_up_slope_drawing_Y	<= '1' when  (oCoord_Y  >= right_up_slope_start_y) and  (oCoord_Y < right_up_slope_end_y) else '0';
	
--	right_up_slope_begin_drawing_X <= '1' when  (oCoord_X  >= (right_up_slope_start_x + right_up_slope_begin_offset)) and  (oCoord_X < (right_up_slope_end_x + right_up_slope_begin_offset)) else '0';
	
	--right_up_slope_drawing_X2	<= '1' when  (oCoord_X  >= right_up_slope_start_x2) and  (oCoord_X < right_up_slope_end_x2) else '0';
   
   tunnel_wall_drawing_X	<= '1' when  (oCoord_X  >= tunnel_wall_start_x) and  (oCoord_X < tunnel_wall_end_x) else '0';
   tunnel_wall_drawing_Y	<= '1' when  (oCoord_Y  >= tunnel_wall_start_y) and  (oCoord_Y < tunnel_wall_end_y) else '0';
   
   stage_left_drawing_X	<= '1' when  (oCoord_X  >= stage_left_start_x) and  (oCoord_X < stage_left_end_x) else '0';
   stage_left_drawing_Y	<= '1' when  (oCoord_Y  >= stage_left_start_y) and  (oCoord_Y < stage_left_end_y) else '0';
   
   stage_right_drawing_X	<= '1' when  (oCoord_X  >= stage_right_start_x) and  (oCoord_X < stage_right_end_x) else '0';
   stage_right_drawing_Y	<= '1' when  (oCoord_Y  >= stage_right_start_y) and  (oCoord_Y < stage_right_end_y) else '0';

	
	start_message_drawing_X	<= '1' when  (oCoord_X  >= start_message_start_x) and  (oCoord_X < start_message_end_x) else '0';
   start_message_drawing_Y	<= '1' when  (oCoord_Y  >= start_message_start_y) and  (oCoord_Y < start_message_end_y) else '0';
	
	game_over_message_drawing_X	<= '1' when  (oCoord_X  >= game_over_message_start_x) and  (oCoord_X < game_over_message_end_x) else '0';
   game_over_message_drawing_Y	<= '1' when  (oCoord_Y  >= game_over_message_start_y) and  (oCoord_Y < game_over_message_end_y) else '0';

	
	
	
	-- calculate offset from start corner 
	left_down_slope_Coord_X 	<= (oCoord_X - left_down_slope_start_x) when ( left_down_slope_drawing_X = '1' and  left_down_slope_drawing_Y = '1'  ) else 0 ; 
	left_down_slope_Coord_Y 	<= (oCoord_Y - left_down_slope_start_y) when ( left_down_slope_drawing_X = '1' and  left_down_slope_drawing_Y = '1'  ) else 0 ;
	
	left_up_slope_Coord_X 	<= (oCoord_X - left_up_slope_start_x) when ( left_up_slope_drawing_X = '1' and  left_up_slope_drawing_Y = '1'  ) else 0 ; 
	left_up_slope_Coord_Y 	<= (oCoord_Y - left_up_slope_start_y) when ( left_up_slope_drawing_X = '1' and  left_up_slope_drawing_Y = '1'  ) else 0 ;
	
	right_down_slope_Coord_X 	<= (oCoord_X - right_down_slope_start_x) when ( right_down_slope_drawing_X = '1' and  right_down_slope_drawing_Y = '1'  ) else 0 ; 
	right_down_slope_Coord_Y 	<= (oCoord_Y - right_down_slope_start_y) when ( right_down_slope_drawing_X = '1' and  right_down_slope_drawing_Y = '1'  ) else 0 ;
	
	right_up_slope_Coord_X 	<= (oCoord_X - right_up_slope_start_x) when ( right_up_slope_drawing_X = '1' and  right_up_slope_drawing_Y = '1'  ) else 0 ; 
	right_up_slope_Coord_Y 	<= (oCoord_Y - right_up_slope_start_y) when ( right_up_slope_drawing_X = '1' and  right_up_slope_drawing_Y = '1'  ) else 0 ;
	
--	right_up_slope_begin_Coord_X <= (oCoord_X - (right_up_slope_start_x + right_up_slope_begin_offset)) when ( right_up_slope_begin_drawing_X = '1' and  right_up_slope_drawing_Y = '1'  ) else 0 ;
--	right_up_slope_Coord_X2 	<= (oCoord_X - right_up_slope_start_x2) when ( right_up_slope_drawing_X2 = '1' and  right_up_slope_drawing_Y = '1'  ) else 0 ; 


	tunnel_wall_Coord_X 	<= (oCoord_X - tunnel_wall_start_x) when ( tunnel_wall_drawing_X = '1' and  tunnel_wall_drawing_Y = '1'  ) else 0 ; 
	tunnel_wall_Coord_Y 	<= (oCoord_Y - tunnel_wall_start_y) when ( tunnel_wall_drawing_X = '1' and  tunnel_wall_drawing_Y = '1'  ) else 0 ;
	
	start_message_Coord_X 	<= (oCoord_X - start_message_start_x) when ( start_message_drawing_X = '1' and  start_message_drawing_Y = '1'  ) else 0 ; 
	start_message_Coord_Y 	<= (oCoord_Y - start_message_start_y) when ( start_message_drawing_X = '1' and  start_message_drawing_Y = '1'  ) else 0 ;
	
	game_over_message_Coord_X 	<= (oCoord_X - game_over_message_start_x) when ( game_over_message_drawing_X = '1' and  game_over_message_drawing_Y = '1'  ) else 0 ; 
	game_over_message_Coord_Y 	<= (oCoord_Y - game_over_message_start_y) when ( game_over_message_drawing_X = '1' and  game_over_message_drawing_Y = '1'  ) else 0 ;
	
	
	-------------------------------------------------------------------
	
	obsticle_up_drawing_X	<= '1' when  (oCoord_X  >= obsticle_up_start_x) and  (oCoord_X < obsticle_up_end_x) else '0';
   obsticle_up_drawing_Y	<= '1' when  (oCoord_Y  >= obsticle_up_start_y) and  (oCoord_Y < obsticle_up_end_y) else '0';

	obsticle_left_up_drawing_X	<= '1' when  (oCoord_X  >= obsticle_left_up_start_x) and  (oCoord_X < obsticle_left_up_end_x) else '0';
   obsticle_left_up_drawing_Y	<= '1' when  (oCoord_Y  >= obsticle_left_up_start_y) and  (oCoord_Y < obsticle_left_up_end_y) else '0';

	obsticle_left_drawing_X	<= '1' when  (oCoord_X  >= obsticle_left_start_x) and  (oCoord_X < obsticle_left_end_x) else '0';
   obsticle_left_drawing_Y	<= '1' when  (oCoord_Y  >= obsticle_left_start_y) and  (oCoord_Y < obsticle_left_end_y) else '0';

	obsticle_left_down_drawing_X	<= '1' when  (oCoord_X  >= obsticle_left_down_start_x) and  (oCoord_X < obsticle_left_down_end_x) else '0';
   obsticle_left_down_drawing_Y	<= '1' when  (oCoord_Y  >= obsticle_left_down_start_y) and  (oCoord_Y < obsticle_left_down_end_y) else '0';

	obsticle_down_drawing_X	<= '1' when  (oCoord_X  >= obsticle_down_start_x) and  (oCoord_X < obsticle_down_end_x) else '0';
   obsticle_down_drawing_Y	<= '1' when  (oCoord_Y  >= obsticle_down_start_y) and  (oCoord_Y < obsticle_down_end_y) else '0';

	obsticle_right_down_drawing_X	<= '1' when  (oCoord_X  >= obsticle_right_down_start_x) and  (oCoord_X < obsticle_right_down_end_x) else '0';
   obsticle_right_down_drawing_Y	<= '1' when  (oCoord_Y  >= obsticle_right_down_start_y) and  (oCoord_Y < obsticle_right_down_end_y) else '0';

	obsticle_right_drawing_X	<= '1' when  (oCoord_X  >= obsticle_right_start_x) and  (oCoord_X < obsticle_right_end_x) else '0';
   obsticle_right_drawing_Y	<= '1' when  (oCoord_Y  >= obsticle_right_start_y) and  (oCoord_Y < obsticle_right_end_y) else '0';

	obsticle_right_up_drawing_X	<= '1' when  (oCoord_X  >= obsticle_right_up_start_x) and  (oCoord_X < obsticle_right_up_end_x) else '0';
   obsticle_right_up_drawing_Y	<= '1' when  (oCoord_Y  >= obsticle_right_up_start_y) and  (oCoord_Y < obsticle_right_up_end_y) else '0';


	-- calculate offset from start corner 
	obsticle_left_up_Coord_X 	<= (oCoord_X - obsticle_left_up_start_x) when ( obsticle_left_up_drawing_X = '1' and  obsticle_left_up_drawing_Y = '1'  ) else 0 ; 
	obsticle_left_up_Coord_Y 	<= (oCoord_Y - obsticle_left_up_start_y) when ( obsticle_left_up_drawing_X = '1' and  obsticle_left_up_drawing_Y = '1'  ) else 0 ;
	
	obsticle_left_down_Coord_X 	<= (oCoord_X - obsticle_left_down_start_x) when ( obsticle_left_down_drawing_X = '1' and  obsticle_left_down_drawing_Y = '1'  ) else 0 ; 
	obsticle_left_down_Coord_Y 	<= (oCoord_Y - obsticle_left_down_start_y) when ( obsticle_left_down_drawing_X = '1' and  obsticle_left_down_drawing_Y = '1'  ) else 0 ;
	
	obsticle_right_down_Coord_X 	<= (oCoord_X - obsticle_right_down_start_x) when ( obsticle_right_down_drawing_X = '1' and  obsticle_right_down_drawing_Y = '1'  ) else 0 ; 
	obsticle_right_down_Coord_Y 	<= (oCoord_Y - obsticle_right_down_start_y) when ( obsticle_right_down_drawing_X = '1' and  obsticle_right_down_drawing_Y = '1'  ) else 0 ;
	
	obsticle_right_up_Coord_X 	<= (oCoord_X - obsticle_right_up_start_x) when ( obsticle_right_up_drawing_X = '1' and  obsticle_right_up_drawing_Y = '1'  ) else 0 ; 
	obsticle_right_up_Coord_Y 	<= (oCoord_Y - obsticle_right_up_start_y) when ( obsticle_right_up_drawing_X = '1' and  obsticle_right_up_drawing_Y = '1'  ) else 0 ;

	
	-------------------------------------------------------------------
	
	-------------------------------------------------------------------
	
	obsticle_2_up_drawing_X	<= '1' when  (oCoord_X  >= obsticle_up_start_x + obsticle_2_x_offset) and  (oCoord_X < obsticle_up_end_x + obsticle_2_x_offset) else '0';
   obsticle_2_up_drawing_Y	<= '1' when  (oCoord_Y  >= obsticle_up_start_y + obsticle_2_y_offset) and  (oCoord_Y < obsticle_up_end_y + obsticle_2_y_offset) else '0';

	obsticle_2_left_up_drawing_X	<= '1' when  (oCoord_X  >= obsticle_left_up_start_x + obsticle_2_x_offset) and  (oCoord_X < obsticle_left_up_end_x + obsticle_2_x_offset) else '0';
   obsticle_2_left_up_drawing_Y	<= '1' when  (oCoord_Y  >= obsticle_left_up_start_y + obsticle_2_y_offset) and  (oCoord_Y < obsticle_left_up_end_y + obsticle_2_y_offset) else '0';

	obsticle_2_left_drawing_X	<= '1' when  (oCoord_X  >= obsticle_left_start_x + obsticle_2_x_offset) and  (oCoord_X < obsticle_left_end_x + obsticle_2_x_offset) else '0';
   obsticle_2_left_drawing_Y	<= '1' when  (oCoord_Y  >= obsticle_left_start_y + obsticle_2_y_offset) and  (oCoord_Y < obsticle_left_end_y + obsticle_2_y_offset) else '0';

	obsticle_2_left_down_drawing_X	<= '1' when  (oCoord_X  >= obsticle_left_down_start_x + obsticle_2_x_offset) and  (oCoord_X < obsticle_left_down_end_x + obsticle_2_x_offset) else '0';
   obsticle_2_left_down_drawing_Y	<= '1' when  (oCoord_Y  >= obsticle_left_down_start_y + obsticle_2_y_offset) and  (oCoord_Y < obsticle_left_down_end_y + obsticle_2_y_offset) else '0';

	obsticle_2_down_drawing_X	<= '1' when  (oCoord_X  >= obsticle_down_start_x + obsticle_2_x_offset) and  (oCoord_X < obsticle_down_end_x + obsticle_2_x_offset) else '0';
   obsticle_2_down_drawing_Y	<= '1' when  (oCoord_Y  >= obsticle_down_start_y + obsticle_2_y_offset) and  (oCoord_Y < obsticle_down_end_y + obsticle_2_y_offset) else '0';

	obsticle_2_right_down_drawing_X	<= '1' when  (oCoord_X  >= obsticle_right_down_start_x + obsticle_2_x_offset) and  (oCoord_X < obsticle_right_down_end_x + obsticle_2_x_offset) else '0';
   obsticle_2_right_down_drawing_Y	<= '1' when  (oCoord_Y  >= obsticle_right_down_start_y + obsticle_2_y_offset) and  (oCoord_Y < obsticle_right_down_end_y + obsticle_2_y_offset) else '0';

	obsticle_2_right_drawing_X	<= '1' when  (oCoord_X  >= obsticle_right_start_x + obsticle_2_x_offset) and  (oCoord_X < obsticle_right_end_x + obsticle_2_x_offset) else '0';
   obsticle_2_right_drawing_Y	<= '1' when  (oCoord_Y  >= obsticle_right_start_y + obsticle_2_y_offset) and  (oCoord_Y < obsticle_right_end_y + obsticle_2_y_offset) else '0';

	obsticle_2_right_up_drawing_X	<= '1' when  (oCoord_X  >= obsticle_right_up_start_x + obsticle_2_x_offset) and  (oCoord_X < obsticle_right_up_end_x + obsticle_2_x_offset) else '0';
   obsticle_2_right_up_drawing_Y	<= '1' when  (oCoord_Y  >= obsticle_right_up_start_y + obsticle_2_y_offset) and  (oCoord_Y < obsticle_right_up_end_y + obsticle_2_y_offset) else '0';


	-- calculate offset from start corner 
	obsticle_2_left_up_Coord_X 	<= (oCoord_X - (obsticle_left_up_start_x + obsticle_2_x_offset)) when ( obsticle_2_left_up_drawing_X = '1' and  obsticle_2_left_up_drawing_Y = '1'  ) else 0 ; 
	obsticle_2_left_up_Coord_Y 	<= (oCoord_Y - (obsticle_left_up_start_y + obsticle_2_y_offset)) when ( obsticle_2_left_up_drawing_X = '1' and  obsticle_2_left_up_drawing_Y = '1'  ) else 0 ;
	
	obsticle_2_left_down_Coord_X 	<= (oCoord_X - (obsticle_left_down_start_x + obsticle_2_x_offset)) when ( obsticle_2_left_down_drawing_X = '1' and  obsticle_2_left_down_drawing_Y = '1'  ) else 0 ; 
	obsticle_2_left_down_Coord_Y 	<= (oCoord_Y - (obsticle_left_down_start_y + obsticle_2_y_offset)) when ( obsticle_2_left_down_drawing_X = '1' and  obsticle_2_left_down_drawing_Y = '1'  ) else 0 ;
	
	obsticle_2_right_down_Coord_X 	<= (oCoord_X - (obsticle_right_down_start_x + obsticle_2_x_offset)) when ( obsticle_2_right_down_drawing_X = '1' and  obsticle_2_right_down_drawing_Y = '1'  ) else 0 ; 
	obsticle_2_right_down_Coord_Y 	<= (oCoord_Y - (obsticle_right_down_start_y + obsticle_2_y_offset)) when ( obsticle_2_right_down_drawing_X = '1' and  obsticle_2_right_down_drawing_Y = '1'  ) else 0 ;
	
	obsticle_2_right_up_Coord_X 	<= (oCoord_X - (obsticle_right_up_start_x + obsticle_2_x_offset)) when ( obsticle_2_right_up_drawing_X = '1' and  obsticle_2_right_up_drawing_Y = '1'  ) else 0 ; 
	obsticle_2_right_up_Coord_Y 	<= (oCoord_Y - (obsticle_right_up_start_y + obsticle_2_y_offset)) when ( obsticle_2_right_up_drawing_X = '1' and  obsticle_2_right_up_drawing_Y = '1'  ) else 0 ;
--------------------------------------------------------------------------------------------------------------------------------------------------------

	--------------------------------------------------------------------------------------------------------------------------------------------------------
	
	obsticle_3_up_drawing_X	<= '1' when  (oCoord_X  >= obsticle_up_start_x + obsticle_3_x_offset) and  (oCoord_X < obsticle_up_end_x + obsticle_3_x_offset) else '0';
   obsticle_3_up_drawing_Y	<= '1' when  (oCoord_Y  >= obsticle_up_start_y + obsticle_3_y_offset) and  (oCoord_Y < obsticle_up_end_y + obsticle_3_y_offset) else '0';

	obsticle_3_left_up_drawing_X	<= '1' when  (oCoord_X  >= obsticle_left_up_start_x + obsticle_3_x_offset) and  (oCoord_X < obsticle_left_up_end_x + obsticle_3_x_offset) else '0';
   obsticle_3_left_up_drawing_Y	<= '1' when  (oCoord_Y  >= obsticle_left_up_start_y + obsticle_3_y_offset) and  (oCoord_Y < obsticle_left_up_end_y + obsticle_3_y_offset) else '0';

	obsticle_3_left_drawing_X	<= '1' when  (oCoord_X  >= obsticle_left_start_x + obsticle_3_x_offset) and  (oCoord_X < obsticle_left_end_x + obsticle_3_x_offset) else '0';
   obsticle_3_left_drawing_Y	<= '1' when  (oCoord_Y  >= obsticle_left_start_y + obsticle_3_y_offset) and  (oCoord_Y < obsticle_left_end_y + obsticle_3_y_offset) else '0';

	obsticle_3_left_down_drawing_X	<= '1' when  (oCoord_X  >= obsticle_left_down_start_x + obsticle_3_x_offset) and  (oCoord_X < obsticle_left_down_end_x + obsticle_3_x_offset) else '0';
   obsticle_3_left_down_drawing_Y	<= '1' when  (oCoord_Y  >= obsticle_left_down_start_y + obsticle_3_y_offset) and  (oCoord_Y < obsticle_left_down_end_y + obsticle_3_y_offset) else '0';

	obsticle_3_down_drawing_X	<= '1' when  (oCoord_X  >= obsticle_down_start_x + obsticle_3_x_offset) and  (oCoord_X < obsticle_down_end_x + obsticle_3_x_offset) else '0';
   obsticle_3_down_drawing_Y	<= '1' when  (oCoord_Y  >= obsticle_down_start_y + obsticle_3_y_offset) and  (oCoord_Y < obsticle_down_end_y + obsticle_3_y_offset) else '0';

	obsticle_3_right_down_drawing_X	<= '1' when  (oCoord_X  >= obsticle_right_down_start_x + obsticle_3_x_offset) and  (oCoord_X < obsticle_right_down_end_x + obsticle_3_x_offset) else '0';
   obsticle_3_right_down_drawing_Y	<= '1' when  (oCoord_Y  >= obsticle_right_down_start_y + obsticle_3_y_offset) and  (oCoord_Y < obsticle_right_down_end_y + obsticle_3_y_offset) else '0';

	obsticle_3_right_drawing_X	<= '1' when  (oCoord_X  >= obsticle_right_start_x + obsticle_3_x_offset) and  (oCoord_X < obsticle_right_end_x + obsticle_3_x_offset) else '0';
   obsticle_3_right_drawing_Y	<= '1' when  (oCoord_Y  >= obsticle_right_start_y + obsticle_3_y_offset) and  (oCoord_Y < obsticle_right_end_y + obsticle_3_y_offset) else '0';

	obsticle_3_right_up_drawing_X	<= '1' when  (oCoord_X  >= obsticle_right_up_start_x + obsticle_3_x_offset) and  (oCoord_X < obsticle_right_up_end_x + obsticle_3_x_offset) else '0';
   obsticle_3_right_up_drawing_Y	<= '1' when  (oCoord_Y  >= obsticle_right_up_start_y + obsticle_3_y_offset) and  (oCoord_Y < obsticle_right_up_end_y + obsticle_3_y_offset) else '0';


	-- calculate offset from start corner 
	obsticle_3_left_up_Coord_X 	<= (oCoord_X - (obsticle_left_up_start_x + obsticle_3_x_offset)) when ( obsticle_3_left_up_drawing_X = '1' and  obsticle_3_left_up_drawing_Y = '1'  ) else 0 ; 
	obsticle_3_left_up_Coord_Y 	<= (oCoord_Y - (obsticle_left_up_start_y + obsticle_3_y_offset)) when ( obsticle_3_left_up_drawing_X = '1' and  obsticle_3_left_up_drawing_Y = '1'  ) else 0 ;
	
	obsticle_3_left_down_Coord_X 	<= (oCoord_X - (obsticle_left_down_start_x + obsticle_3_x_offset)) when ( obsticle_3_left_down_drawing_X = '1' and  obsticle_3_left_down_drawing_Y = '1'  ) else 0 ; 
	obsticle_3_left_down_Coord_Y 	<= (oCoord_Y - (obsticle_left_down_start_y + obsticle_3_y_offset)) when ( obsticle_3_left_down_drawing_X = '1' and  obsticle_3_left_down_drawing_Y = '1'  ) else 0 ;
	
	obsticle_3_right_down_Coord_X 	<= (oCoord_X - (obsticle_right_down_start_x + obsticle_3_x_offset)) when ( obsticle_3_right_down_drawing_X = '1' and  obsticle_3_right_down_drawing_Y = '1'  ) else 0 ; 
	obsticle_3_right_down_Coord_Y 	<= (oCoord_Y - (obsticle_right_down_start_y + obsticle_3_y_offset)) when ( obsticle_3_right_down_drawing_X = '1' and  obsticle_3_right_down_drawing_Y = '1'  ) else 0 ;
	
	obsticle_3_right_up_Coord_X 	<= (oCoord_X - (obsticle_right_up_start_x + obsticle_3_x_offset)) when ( obsticle_3_right_up_drawing_X = '1' and  obsticle_3_right_up_drawing_Y = '1'  ) else 0 ; 
	obsticle_3_right_up_Coord_Y 	<= (oCoord_Y - (obsticle_right_up_start_y + obsticle_3_y_offset)) when ( obsticle_3_right_up_drawing_X = '1' and  obsticle_3_right_up_drawing_Y = '1'  ) else 0 ;

	
	-------------------------------------------------------------------


	
process ( RESETn, CLK)

  		
   begin
		
	if RESETn = '0' then
	    mVGA_RGB	<=  (others => '0') ; 	
		 drawing_request	<=  '0' ;
		 sigSpaceWasPressed <= '0';
		 sigGameOver <= '0';

	elsif rising_edge(CLK) then
	
		sig_draw_req <= '0';
		sig_bounce_type <= no_bounce;
		
		if (space_was_pressed = '1') then
			sigSpaceWasPressed <= '1';
		end if;
		
		if (game_over = '1') then
			sigGameOver <= '1';
		end if;
		

		
		if ( (floor_drawing_X ='1') and (floor_drawing_Y = '1') ) then
			sig_draw_req <= '1';
			sig_draw_data <= floor_color;
			if (oCoord_Y <= fell_to_pit_upper_Y_bound) then
				sig_bounce_type <= floor_bounce_type;
			else
				sig_bounce_type <= death;
			end if;
			
		end if;
		

		if ((ceiling_drawing_X ='1') and (ceiling_drawing_Y = '1') ) then
			sig_draw_req <= '1';
			sig_draw_data <= ceiling_color;
			sig_bounce_type <= ceiling_bounce_type;
		end if;	
		

		if ((left_wall_drawing_X ='1') and (left_wall_drawing_Y = '1')) then
			sig_draw_req <= '1';
			sig_draw_data <= left_wall_color;
			sig_bounce_type <= left_wall_bounce_type;
		end if;

		if ((right_wall_drawing_X ='1') and (right_wall_drawing_Y = '1')) then
			sig_draw_req <= '1';
			sig_draw_data <= right_wall_color;
			sig_bounce_type <= right_wall_bounce_type;
		end if;
		
		if ( (stage_left_drawing_X ='1') and (stage_left_drawing_Y = '1') ) then
			sig_draw_req <= '1';
			sig_draw_data <= stage_left_color;
			if fell_to_pit = '1' then
				sig_bounce_type <= stage_left_bounce_type2;
			else
				sig_bounce_type <= stage_left_bounce_type1;
			end if;
		end if;
		
		if ( (stage_right_drawing_X ='1') and (stage_right_drawing_Y = '1') ) then
			sig_draw_req <= '1';
			sig_draw_data <= stage_right_color;
			if fell_to_pit = '1' then
				sig_bounce_type <= stage_right_bounce_type2;
			else
				sig_bounce_type <= stage_right_bounce_type1;
			end if;
		end if;
		
		----------------------------------------------------------------------------
		
		if ((left_down_slope_drawing_X ='1') and (left_down_slope_drawing_Y = '1')) then
			sig_draw_req <= left_down_slope_object(left_down_slope_Coord_Y,left_down_slope_Coord_X);
			sig_draw_data <= left_down_slope_color;
			if left_down_slope_object(left_down_slope_Coord_Y,left_down_slope_Coord_X) = '1' then
				sig_bounce_type <= left_down_slope_bounce_type;
			else
				sig_bounce_type <= no_bounce;
			end if;
		end if;
		
		if ((left_up_slope_drawing_X ='1') and (left_up_slope_drawing_Y = '1')) then
			sig_draw_req <= left_up_slope_object(left_up_slope_Coord_Y,left_up_slope_Coord_X);
			sig_draw_data <= left_up_slope_color;
			if left_up_slope_object(left_up_slope_Coord_Y,left_up_slope_Coord_X) = '1' then
				sig_bounce_type <= left_up_slope_bounce_type;
			else
				sig_bounce_type <= no_bounce;
			end if;
		end if;
		
		if ((right_down_slope_drawing_X ='1') and (right_down_slope_drawing_Y = '1')) then
			sig_draw_req <= right_down_slope_object(right_down_slope_Coord_Y, right_down_slope_Coord_X);
			sig_draw_data <= right_down_slope_color;
			if right_down_slope_object(right_down_slope_Coord_Y, right_down_slope_Coord_X) = '1' then
				sig_bounce_type <= right_down_slope_bounce_type;
			else
				sig_bounce_type <= no_bounce;
			end if;
		end if;
		
		
		--if ((right_up_slope_drawing_X ='1' or right_up_slope_drawing_X2 = '1') and (right_up_slope_drawing_Y = '1')) then
		--	sig_draw_data <= right_up_slope_color;
		--	if (game_started = '0') then
		--		sig_draw_req <= right_up_slope_object(right_up_slope_Coord_Y,right_up_slope_Coord_X);
		--		if right_up_slope_object(right_up_slope_Coord_Y,right_up_slope_Coord_X) = '1' then
		--			sig_bounce_type <= right_up_slope_bounce_type;
		--		else
		--			sig_bounce_type <= no_bounce;
		--		end if;
		--	else
		--		sig_draw_req <= right_up_slope_object(right_up_slope_Coord_Y,right_up_slope_Coord_X2);
		--		if right_up_slope_object(right_up_slope_Coord_Y,right_up_slope_Coord_X2) = '1' then
		--			sig_bounce_type <= right_up_slope_bounce_type;
		--		else
		--			sig_bounce_type <= no_bounce;
		--		end if;
		--
		--	end if;
		--end if;
		
--		if (game_started = '0') then
			if ((right_up_slope_drawing_X ='1' ) and (right_up_slope_drawing_Y = '1')) then
				sig_draw_req <= right_up_slope_object(right_up_slope_Coord_Y,right_up_slope_Coord_X);
				sig_draw_data <= right_up_slope_color;
				if right_up_slope_object(right_up_slope_Coord_Y,right_up_slope_Coord_X) = '1' then
					sig_bounce_type <= right_up_slope_bounce_type;
				else
					sig_bounce_type <= no_bounce;
				end if;
			end if;
--		else
--			if ((right_up_slope_begin_drawing_X ='1' ) and (right_up_slope_drawing_Y = '1')) then
--				sig_draw_req <= right_up_slope_object(right_up_slope_Coord_Y,right_up_slope_begin_Coord_X);
--				sig_draw_data <= right_up_slope_color;
--				if right_up_slope_object(right_up_slope_Coord_Y,right_up_slope_begin_Coord_X) = '1' then
--					sig_bounce_type <= left_up_slope_bounce_type;
--				else
--					sig_bounce_type <= no_bounce;
--				end if;
--			end if;
--		end if;
			

		
		
		if ((tunnel_wall_drawing_X ='1') and (tunnel_wall_drawing_Y = '1')) then
			if game_started = '1' then 
				sig_draw_req <= '1';
				sig_bounce_type <= tunnel_wall_bounce_type;
			else
				sig_draw_req <= tunnel_wall_object(tunnel_wall_Coord_Y,tunnel_wall_Coord_X);
				if tunnel_wall_object(tunnel_wall_Coord_Y,tunnel_wall_Coord_X) = '1' then
					sig_bounce_type <= tunnel_wall_bounce_type;
				else
					sig_bounce_type <= no_bounce;
				end if;
			end if;
			sig_draw_data <= tunnel_wall_color;
		end if;

		----------------------------------------------------------------------------
		if ((obsticle_up_drawing_X ='1') and (obsticle_up_drawing_Y = '1')) then			-- obsticle up
			sig_draw_req <= '1';
			sig_draw_data <= obsticle_up_color;
			sig_bounce_type <= obsticle_up_bounce_type;
		end if;

		if ((obsticle_left_up_drawing_X ='1') and (obsticle_left_up_drawing_Y = '1')) then			-- obsticle left up
			sig_draw_req <= obsticle_left_up_mask(obsticle_left_up_Coord_Y,obsticle_left_up_Coord_X);
			sig_draw_data <= obsticle_left_up_color;
			if obsticle_left_up_mask(obsticle_left_up_Coord_Y,obsticle_left_up_Coord_X) = '1' then
				sig_bounce_type <= obsticle_left_up_bounce_type;
			else
				sig_bounce_type <= no_bounce;
			end if;
		end if;

		if ((obsticle_left_drawing_X ='1') and (obsticle_left_drawing_Y = '1')) then		-- obsticke left
			sig_draw_req <= '1';
			sig_draw_data <= obsticle_left_color;
			sig_bounce_type <= obsticle_left_bounce_type;
		end if;

		if ((obsticle_left_down_drawing_X ='1') and (obsticle_left_down_drawing_Y = '1')) then			-- obsticle left down
			sig_draw_req <= obsticle_left_down_mask(obsticle_left_down_Coord_Y,obsticle_left_down_Coord_X);
			sig_draw_data <= obsticle_left_down_color;
			if obsticle_left_down_mask(obsticle_left_down_Coord_Y,obsticle_left_down_Coord_X) = '1' then
				sig_bounce_type <= obsticle_left_down_bounce_type;
			else
				sig_bounce_type <= no_bounce;
			end if;
		end if;

		if ((obsticle_down_drawing_X ='1') and (obsticle_down_drawing_Y = '1')) then		-- obsticle down
			sig_draw_req <= '1';
			sig_draw_data <= obsticle_down_color;
			sig_bounce_type <= obsticle_down_bounce_type;
		end if;

		if ((obsticle_right_down_drawing_X ='1') and (obsticle_right_down_drawing_Y = '1')) then			-- obsticle right down
			sig_draw_req <= obsticle_right_down_mask(obsticle_right_down_Coord_Y,obsticle_right_down_Coord_X);
			sig_draw_data <= obsticle_right_down_color;
			if obsticle_right_down_mask(obsticle_right_down_Coord_Y,obsticle_right_down_Coord_X) = '1' then
				sig_bounce_type <= obsticle_right_down_bounce_type;
			else
				sig_bounce_type <= no_bounce;
			end if;
		end if;

		if ((obsticle_right_drawing_X ='1') and (obsticle_right_drawing_Y = '1')) then		-- obsticle right
			sig_draw_req <= '1';
			sig_draw_data <= obsticle_right_color;
			sig_bounce_type <= obsticle_right_bounce_type;
		end if;

		if ((obsticle_right_up_drawing_X ='1') and (obsticle_right_up_drawing_Y = '1')) then		-- obsticle right up
			sig_draw_req <= obsticle_right_up_mask(obsticle_right_up_Coord_Y,obsticle_right_up_Coord_X);
			sig_draw_data <= obsticle_right_up_color;
			if obsticle_right_up_mask(obsticle_right_up_Coord_Y,obsticle_right_up_Coord_X) = '1' then
				sig_bounce_type <= obsticle_right_up_bounce_type;
			else
				sig_bounce_type <= no_bounce;
			end if;
		end if;
		
		-----------------------------------------------------------------------------
		
		----------------------------------------------------------------------------
		if ((obsticle_2_up_drawing_X ='1') and (obsticle_2_up_drawing_Y = '1')) then			-- obsticle up
			sig_draw_req <= '1';
			sig_draw_data <= obsticle_up_color;
			sig_bounce_type <= obsticle_up_bounce_type;
		end if;

		if ((obsticle_2_left_up_drawing_X ='1') and (obsticle_2_left_up_drawing_Y = '1')) then			-- obsticle left up
			sig_draw_req <= obsticle_left_up_mask(obsticle_2_left_up_Coord_Y,obsticle_2_left_up_Coord_X);
			sig_draw_data <= obsticle_left_up_color;
			if obsticle_left_up_mask(obsticle_2_left_up_Coord_Y,obsticle_2_left_up_Coord_X) = '1' then
				sig_bounce_type <= obsticle_left_up_bounce_type;
			else
				sig_bounce_type <= no_bounce;
			end if;
		end if;

		if ((obsticle_2_left_drawing_X ='1') and (obsticle_2_left_drawing_Y = '1')) then		-- obsticke left
			sig_draw_req <= '1';
			sig_draw_data <= obsticle_left_color;
			sig_bounce_type <= obsticle_left_bounce_type;
		end if;

		if ((obsticle_2_left_down_drawing_X ='1') and (obsticle_2_left_down_drawing_Y = '1')) then			-- obsticle left down
			sig_draw_req <= obsticle_left_down_mask(obsticle_2_left_down_Coord_Y,obsticle_2_left_down_Coord_X);
			sig_draw_data <= obsticle_left_down_color;
			if obsticle_left_down_mask(obsticle_2_left_down_Coord_Y,obsticle_2_left_down_Coord_X) = '1' then
				sig_bounce_type <= obsticle_left_down_bounce_type;
			else
				sig_bounce_type <= no_bounce;
			end if;
		end if;

		if ((obsticle_2_down_drawing_X ='1') and (obsticle_2_down_drawing_Y = '1')) then		-- obsticle down
			sig_draw_req <= '1';
			sig_draw_data <= obsticle_down_color;
			sig_bounce_type <= obsticle_down_bounce_type;
		end if;

		if ((obsticle_2_right_down_drawing_X ='1') and (obsticle_2_right_down_drawing_Y = '1')) then			-- obsticle right down
			sig_draw_req <= obsticle_right_down_mask(obsticle_2_right_down_Coord_Y,obsticle_2_right_down_Coord_X);
			sig_draw_data <= obsticle_right_down_color;
			if obsticle_right_down_mask(obsticle_2_right_down_Coord_Y,obsticle_2_right_down_Coord_X) = '1' then
				sig_bounce_type <= obsticle_right_down_bounce_type;
			else
				sig_bounce_type <= no_bounce;
			end if;
		end if;

		if ((obsticle_2_right_drawing_X ='1') and (obsticle_2_right_drawing_Y = '1')) then		-- obsticle right
			sig_draw_req <= '1';
			sig_draw_data <= obsticle_right_color;
			sig_bounce_type <= obsticle_right_bounce_type;
		end if;

		if ((obsticle_2_right_up_drawing_X ='1') and (obsticle_2_right_up_drawing_Y = '1')) then		-- obsticle right up
			sig_draw_req <= obsticle_right_up_mask(obsticle_2_right_up_Coord_Y,obsticle_2_right_up_Coord_X);
			sig_draw_data <= obsticle_right_up_color;
			if obsticle_right_up_mask(obsticle_2_right_up_Coord_Y,obsticle_2_right_up_Coord_X) = '1' then
				sig_bounce_type <= obsticle_right_up_bounce_type;
			else
				sig_bounce_type <= no_bounce;
			end if;
		end if;
		
		----------------------------------------------------------------------------------------------
				----------------------------------------------------------------------------
		if ((obsticle_3_up_drawing_X ='1') and (obsticle_3_up_drawing_Y = '1')) then			-- obsticle up
			sig_draw_req <= '1';
			sig_draw_data <= obsticle_up_color;
			sig_bounce_type <= obsticle_up_bounce_type;
		end if;

		if ((obsticle_3_left_up_drawing_X ='1') and (obsticle_3_left_up_drawing_Y = '1')) then			-- obsticle left up
			sig_draw_req <= obsticle_left_up_mask(obsticle_3_left_up_Coord_Y,obsticle_3_left_up_Coord_X);
			sig_draw_data <= obsticle_left_up_color;
			if obsticle_left_up_mask(obsticle_3_left_up_Coord_Y,obsticle_3_left_up_Coord_X) = '1' then
				sig_bounce_type <= obsticle_left_up_bounce_type;
			else
				sig_bounce_type <= no_bounce;
			end if;
		end if;

		if ((obsticle_3_left_drawing_X ='1') and (obsticle_3_left_drawing_Y = '1')) then		-- obsticke left
			sig_draw_req <= '1';
			sig_draw_data <= obsticle_left_color;
			sig_bounce_type <= obsticle_left_bounce_type;
		end if;

		if ((obsticle_3_left_down_drawing_X ='1') and (obsticle_3_left_down_drawing_Y = '1')) then			-- obsticle left down
			sig_draw_req <= obsticle_left_down_mask(obsticle_3_left_down_Coord_Y,obsticle_3_left_down_Coord_X);
			sig_draw_data <= obsticle_left_down_color;
			if obsticle_left_down_mask(obsticle_3_left_down_Coord_Y,obsticle_3_left_down_Coord_X) = '1' then
				sig_bounce_type <= obsticle_left_down_bounce_type;
			else
				sig_bounce_type <= no_bounce;
			end if;
		end if;

		if ((obsticle_3_down_drawing_X ='1') and (obsticle_3_down_drawing_Y = '1')) then		-- obsticle down
			sig_draw_req <= '1';
			sig_draw_data <= obsticle_down_color;
			sig_bounce_type <= obsticle_down_bounce_type;
		end if;

		if ((obsticle_3_right_down_drawing_X ='1') and (obsticle_3_right_down_drawing_Y = '1')) then			-- obsticle right down
			sig_draw_req <= obsticle_right_down_mask(obsticle_3_right_down_Coord_Y,obsticle_3_right_down_Coord_X);
			sig_draw_data <= obsticle_right_down_color;
			if obsticle_right_down_mask(obsticle_3_right_down_Coord_Y,obsticle_3_right_down_Coord_X) = '1' then
				sig_bounce_type <= obsticle_right_down_bounce_type;
			else
				sig_bounce_type <= no_bounce;
			end if;
		end if;

		if ((obsticle_3_right_drawing_X ='1') and (obsticle_3_right_drawing_Y = '1')) then		-- obsticle right
			sig_draw_req <= '1';
			sig_draw_data <= obsticle_right_color;
			sig_bounce_type <= obsticle_right_bounce_type;
		end if;

		if ((obsticle_3_right_up_drawing_X ='1') and (obsticle_3_right_up_drawing_Y = '1')) then		-- obsticle right up
			sig_draw_req <= obsticle_right_up_mask(obsticle_3_right_up_Coord_Y,obsticle_3_right_up_Coord_X);
			sig_draw_data <= obsticle_right_up_color;
			if obsticle_right_up_mask(obsticle_3_right_up_Coord_Y,obsticle_3_right_up_Coord_X) = '1' then
				sig_bounce_type <= obsticle_right_up_bounce_type;
			else
				sig_bounce_type <= no_bounce;
			end if;
		end if;

		--------------------------------------------------------------------------------------------------------------------
		
		
		if ( (sigSpaceWasPressed = '0') and (start_message_drawing_X = '1') and (start_message_drawing_Y = '1') ) then
			sig_draw_req <= start_message_object(start_message_Coord_Y,start_message_Coord_X);
			sig_draw_data <= start_message_color;
			sig_bounce_type <= start_message_bounce_type;
		end if;
		
		if ( (sigGameOver = '1') and (game_over_message_drawing_X = '1') and (game_over_message_drawing_Y = '1') ) then
			sig_draw_req <= game_over_message_object(start_message_Coord_Y,start_message_Coord_X);
			sig_draw_data <= game_over_message_color;
			sig_bounce_type <= game_over_message_bounce_type;
		end if;
		
		-----------------------------------------------------------------------------

	
			mVGA_RGB	<=  sig_draw_data;	--get from colors table 
			drawing_request	<=  sig_draw_req ; -- get from mask table if inside rectangle
			bounce_type <= sig_bounce_type;
	end if;

  end process;

		
end architecture;	