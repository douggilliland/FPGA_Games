library verilog;
use verilog.vl_types.all;
entity PushBox_vlg_vec_tst is
end PushBox_vlg_vec_tst;
