----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    09:01:08 05/25/2015 
-- Design Name: 
-- Module Name:    Rom_laser_text - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Rom_laser_text is
 Port ( Hposition   : in  STD_LOGIC_VECTOR(10 downto 0);
		  Vposition   : in  STD_LOGIC_VECTOR(9 downto 0);
		  VIDON       : in  STD_LOGIC;
		  enable_game : in  STD_LOGIC;
        obj_rgb     : out  STD_LOGIC;
		  obj_on      : out  STD_LOGIC );
end Rom_laser_text;

architecture Behavioral of Rom_laser_text is

type ROM is array(0 to 39) of std_logic_vector(99 downto 0);
constant content : ROM := (

0 =>"1111110000000000000000000001111000000000001111111111111111001111111111111111110011111110000000000000",
1 =>"1111110000000000000000000011111100000000011111111111111111001111111111111111110011111111100000000000",
2 =>"1111110000000000000000000111111110000000111111111111111111001111111111111111110011111111111000000000",
3 =>"1111110000000000000000000111111110000000111111111111111111001111111111111111110011111111111000000000",
4 =>"1111110000000000000000000111111110000000111111100000000000001111110000000000000011111111111110000000",
5 =>"1111110000000000000000000111111110000000111111000000000000001111110000000000000011111111111111000000",
6 =>"1111110000000000000000001111111111000000111111000000000000001111110000000000000011111100000011110000",
7 =>"1111110000000000000000001111111111000000111111000000000000001111110000000000000011111100000011111000",
8 =>"1111110000000000000000001111111111100000111111000000000000001111110000000000000011111100000001111110",
9 =>"1111110000000000000000111111111111110000111111000000000000001111110000000000000011111100000000111110",
10=>"1111110000000000000000111111001111110000111111000000000000001111110000000000000011111100000000011111",
11=>"1111110000000000000000111111001111110000111111000000000000001111110000000000000011111100000000011111",
12=>"1111110000000000000001111110000111111000011111100000000000001111110000000000000011111100000000011111",
13=>"1111110000000000000001111110000111111000001111110000000000001111110000000000000011111100000000111110",
14=>"1111110000000000000001111110000111111000000011111100000000001111110000000000000011111100000001111100",
15=>"1111110000000000000011111110000111111100000011111100000000001111110000000000000011111100000001111100",
16=>"1111110000000000000011111110000111111100000001111110000000001111110000000000000011111100000011111000",
17=>"1111110000000000000011111111111111111100000001111110000000001111111111111100000011111100000111110000",
18=>"1111110000000000000011111111111111111100000000111111000000001111111111111100000011111100011111000000",
19=>"1111110000000000000011111111111111111100000000111111000000001111111111111100000011111100111110000000",
20=>"1111110000000000000011111111111111111100000000011111100000001111111111111100000011111101111100000000",
21=>"1111110000000000000011111110000111111100000000011111100000001111110000000000000011111111111000000000",
22=>"1111110000000000000011111110000111111100000000001111110000001111110000000000000011111111111000000000",
23=>"1111110000000000000011111110000111111100000000001111110000001111110000000000000011111111111000000000",
24=>"1111110000000000000011111110000111111100000000000111111000001111110000000000000011111111111000000000",
25=>"1111110000000000000011111110000111111100000000000111111000001111110000000000000011111101111100000000",
26=>"1111110000000000000011111110000111111100000000000011111100001111110000000000000011111101111100000000",
27=>"1111110000000000000011111110000111111100000000000011111100001111110000000000000011111100111110000000",
28=>"1111110000000000000011111110000111111100000000000001111110001111110000000000000011111100111110000000",
29=>"1111110000000000000011111110000111111100000000000000111111001111110000000000000011111100011111000000",
30=>"1111110000000000000011111110000111111100000000000000111111001111110000000000000011111100011111000000",
31=>"1111110000000000000011111110000111111100000000000000111111001111110000000000000011111100001111100000",
32=>"1111110000000000000011111110000111111100000000000000111111001111110000000000000011111100001111100000",
33=>"1111110000000000000011111110000111111100000000000000111111001111110000000000000011111100000111111000",
34=>"1111110000000000000011111110000111111100000000000000111111001111110000000000000011111100000111111000",
35=>"1111110000000000000011111110000111111100000000000000111111001111110000000000000011111100000011111100",
36=>"1111110000000000000011111110000111111100000000000001111111001111110000000000000011111100000011111100",
37=>"1111111111111111110011111110000111111100111111111111111111001111111111111111110011111100000001111110",
38=>"1111111111111111110011111110000111111100111111111111111111001111111111111111110011111100000001111110",
39=>"1111111111111111110011111110000111111100111111111111111110001111111111111111110011111100000000111111"

);

signal data_line : std_logic_vector(0 to 99);
constant Hstart : std_logic_vector(10 downto 0) := "10001001100"; -- 1100
constant Hend : std_logic_vector(10 downto 0)   := "10010110000"; -- 1200
constant Vstart : std_logic_vector(9 downto 0)  := "0000110010"; -- 50
constant Vend :std_logic_vector(9 downto 0)     := "0001011010"; -- 90

signal obj_row :  STD_LOGIC_VECTOR (10 downto 0);
signal obj_col :  STD_LOGIC_VECTOR (9 downto 0);

signal obj_on_sig : std_logic := '0';
signal object_rgb : std_logic := '0';

begin

process(VIDON, enable_game, Hposition, Vposition)

begin

    object_rgb <= '0';
	 obj_on_sig <= '0';
	 
	 if VIDON = '1' and enable_game = '1' then
	     	  if (Hposition >= Hstart and Hposition < Hend) and
	           (Vposition >= Vstart  and Vposition < Vend) then
		  
					  obj_on_sig <= '1';
					  obj_row <= (Hposition - Hstart);
					  obj_col <= (Vposition - Vstart);
					  
					  data_line <= content(conv_integer(obj_col));
		  
		           object_rgb <= data_line(conv_integer(obj_row));
					  
	        end if;
   
	  end if;

end process;
obj_rgb <= object_rgb;
obj_on <= obj_on_sig;

end Behavioral;
