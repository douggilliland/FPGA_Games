library IEEE;
use IEEE.STD_LOGIC_1164.all;
entity logo2 is
port 	(
		
	   CLK  		: in std_logic;
		RESETn		: in std_logic;
		oCoord_X	: in integer;
		oCoord_Y	: in integer;
		ObjectStartX	: in integer;
		ObjectStartY 	: in integer;
		drawing_request	: out std_logic ;
		mVGA_RGB 	: out std_logic_vector(7 downto 0) 
	);
end entity;


architecture behav of logo2 is 

constant object_X_size : integer := 544;
constant object_Y_size : integer := 219;
type ram_array is array(0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic_vector(7 downto 0);
constant object_colors: ram_array := (
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"b6",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b7",x"b7",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"6d",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"24",x"24",x"49",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"96",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"24",x"00",x"00",x"24",x"24",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"91",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"49",x"24",x"00",x"00",x"24",x"00",x"00",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"49",x"4d",x"6d",x"6d",x"6d",x"6d",x"91",x"92",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"49",x"24",x"00",x"24",x"49",x"6d",x"24",x"00",x"24",x"49",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"49",x"24",x"00",x"00",x"6d",x"b6",x"db",x"49",x"00",x"00",x"24",x"49",x"6d",x"6d",x"6d",x"92",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"6d",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"92",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"24",x"00",x"00",x"00",x"24",x"b6",x"ff",x"ff",x"92",x"24",x"00",x"00",x"49",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"48",x"49",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"92",x"db",x"ff",x"ff",x"b6",x"49",x"00",x"00",x"24",x"49",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"48",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"49",x"db",x"ff",x"ff",x"ff",x"db",x"6d",x"00",x"00",x"24",x"24",x"49",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"92",x"92",x"92",x"6d",x"49",x"24",x"00",x"00",x"00",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"48",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"da",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"49",x"b2",x"ff",x"ff",x"ff",x"ff",x"ff",x"b6",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"24",x"00",x"00",x"00",x"49",x"4a",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"8d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"ba",x"ba",x"ba",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"bb",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"b7",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b7",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"96",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"4d",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"92",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"24",x"00",x"00",x"24",x"24",x"49",x"49",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"bb",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"bb",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"49",x"49",x"24",x"00",x"00",x"25",x"72",x"db",x"92",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"45",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"71",x"71",x"71",x"91",x"91",x"91",x"91",x"91",x"91",x"91",x"92",x"92",x"92",x"92",x"92",x"92",x"71",x"71",x"71",x"72",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"96",x"b6",x"96",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b7",x"d7",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"b6",x"92",x"b6",x"b6",x"92",x"92",x"92",x"92",x"6d",x"72",x"92",x"92",x"92",x"96",x"96",x"96",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b7",x"b7",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"96",x"71",x"6d",x"6d",x"6d",x"6d",x"69",x"69",x"69",x"49",x"49",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"04",x"72",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"6d",x"20",x"00",x"00",x"24",x"24",x"49",x"49",x"6d",x"6d",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"d7",x"b7",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b7",x"b7",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b7",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b7",x"b7",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"92",x"6d",x"6d",x"49",x"49",x"24",x"00",x"00",x"25",x"92",x"ff",x"db",x"72",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"25",x"45",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"96",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b7",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"4d",x"4d",x"49",x"49",x"49",x"49",x"49",x"44",x"24",x"29",x"28",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"49",x"b6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"b6",x"49",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"b2",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"92",x"6d",x"6d",x"49",x"24",x"24",x"00",x"00",x"49",x"b7",x"ff",x"ff",x"db",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"45",x"45",x"45",x"49",x"49",x"49",x"69",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"69",x"69",x"69",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"72",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"91",x"71",x"6d",x"92",x"92",x"92",x"6e",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6e",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"49",x"49",x"6d",x"6d",x"71",x"92",x"92",x"96",x"96",x"b6",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6e",x"6d",x"6d",x"6d",x"6e",x"6e",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"6d",x"69",x"49",x"49",x"29",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"72",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"6d",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6e",x"6e",x"6e",x"6e",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"72",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"92",x"6d",x"6d",x"49",x"24",x"00",x"00",x"00",x"49",x"db",x"ff",x"ff",x"ff",x"b2",x"69",x"45",x"00",x"00",x"00",x"00",x"04",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"45",x"49",x"49",x"45",x"45",x"45",x"45",x"45",x"45",x"49",x"49",x"49",x"48",x"48",x"48",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"48",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6e",x"8e",x"8e",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"44",x"49",x"49",x"6d",x"92",x"92",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"92",x"91",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"6d",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"92",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"91",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"91",x"92",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"71",x"91",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"24",x"00",x"00",x"00",x"49",x"d7",x"ff",x"ff",x"ff",x"fa",x"d6",x"92",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"69",x"69",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"44",x"49",x"69",x"6d",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b7",x"b6",x"b6",x"92",x"92",x"91",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"4d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"44",x"49",x"44",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"96",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"b6",x"49",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"b6",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"4d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"24",x"00",x"00",x"00",x"49",x"b7",x"ff",x"ff",x"fa",x"fa",x"fa",x"d6",x"b2",x"49",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"04",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"49",x"24",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"24",x"44",x"49",x"69",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b7",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"25",x"49",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"29",x"48",x"48",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"00",x"00",x"00",x"20",x"44",x"89",x"b2",x"92",x"6d",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"48",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"48",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"24",x"00",x"00",x"00",x"25",x"92",x"ff",x"ff",x"fa",x"d5",x"d5",x"fa",x"fb",x"d6",x"92",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"00",x"00",x"92",x"b6",x"92",x"00",x"00",x"00",x"24",x"44",x"49",x"49",x"49",x"6d",x"6d",x"71",x"72",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"d7",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"04",x"00",x"00",x"20",x"40",x"84",x"a9",x"f6",x"fb",x"ff",x"ff",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"48",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"92",x"6d",x"6d",x"49",x"24",x"00",x"00",x"00",x"00",x"6e",x"ff",x"ff",x"fa",x"b1",x"b1",x"d5",x"fa",x"fb",x"db",x"b6",x"8e",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"25",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"24",x"db",x"ff",x"db",x"24",x"00",x"00",x"00",x"24",x"24",x"44",x"49",x"49",x"49",x"6d",x"6d",x"72",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b7",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"25",x"49",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"24",x"04",x"00",x"00",x"40",x"60",x"a0",x"c5",x"ee",x"f7",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"6d",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"92",x"6d",x"6d",x"49",x"24",x"24",x"00",x"00",x"00",x"45",x"db",x"ff",x"ff",x"d5",x"b1",x"b1",x"f5",x"fa",x"ff",x"fb",x"f7",x"b2",x"8e",x"69",x"25",x"25",x"20",x"00",x"00",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"20",x"20",x"24",x"24",x"25",x"25",x"25",x"25",x"25",x"49",x"6d",x"6d",x"6e",x"8e",x"92",x"92",x"8e",x"6e",x"69",x"49",x"45",x"25",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"49",x"ff",x"ff",x"ff",x"4d",x"04",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"49",x"4d",x"6d",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"24",x"04",x"00",x"00",x"20",x"60",x"a0",x"c0",x"c4",x"e5",x"ed",x"f6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"b6",x"92",x"6d",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"92",x"db",x"ff",x"fb",x"d5",x"b0",x"b0",x"d1",x"f5",x"f6",x"fa",x"fb",x"fb",x"fb",x"fb",x"d7",x"b6",x"92",x"92",x"8e",x"8e",x"8e",x"92",x"92",x"92",x"b2",x"b2",x"b6",x"d6",x"d6",x"fb",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"db",x"b6",x"92",x"6d",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"25",x"25",x"25",x"45",x"45",x"25",x"25",x"25",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"49",x"b6",x"ff",x"ff",x"ff",x"96",x"4d",x"04",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"49",x"49",x"49",x"69",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"49",x"6d",x"6d",x"91",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"40",x"80",x"c4",x"e5",x"e0",x"c0",x"c4",x"c9",x"f2",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"92",x"6d",x"6d",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"25",x"45",x"45",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"25",x"25",x"25",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"92",x"92",x"6d",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"6e",x"b7",x"ff",x"ff",x"fa",x"d5",x"b0",x"d0",x"d0",x"f1",x"f5",x"fa",x"fa",x"fa",x"ff",x"ff",x"fb",x"db",x"db",x"da",x"da",x"db",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"ff",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"db",x"b6",x"92",x"6d",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"49",x"6e",x"6e",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b7",x"b7",x"b6",x"b6",x"b6",x"92",x"92",x"6e",x"6e",x"6e",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"92",x"ff",x"ff",x"ff",x"ff",x"df",x"96",x"29",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"49",x"6d",x"6e",x"6e",x"6e",x"92",x"92",x"92",x"92",x"92",x"6e",x"6e",x"6e",x"8e",x"8e",x"8e",x"8e",x"8e",x"8e",x"8e",x"8e",x"8e",x"8e",x"8e",x"8e",x"92",x"6e",x"6e",x"49",x"25",x"00",x"00",x"00",x"24",x"49",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"24",x"24",x"24",x"00",x"00",x"20",x"40",x"a4",x"c4",x"e4",x"e0",x"e0",x"c0",x"c5",x"c9",x"f6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"92",x"6d",x"6d",x"49",x"49",x"00",x"00",x"24",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"49",x"49",x"6e",x"8e",x"92",x"92",x"92",x"92",x"b2",x"92",x"92",x"92",x"6e",x"6e",x"6d",x"49",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"49",x"6d",x"6e",x"92",x"92",x"92",x"92",x"96",x"92",x"92",x"92",x"92",x"6e",x"6e",x"49",x"49",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"24",x"00",x"00",x"00",x"00",x"25",x"92",x"fb",x"ff",x"fb",x"f9",x"b0",x"ac",x"cc",x"d0",x"f0",x"f4",x"f5",x"f5",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fe",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f5",x"d5",x"d5",x"d5",x"d5",x"d5",x"d5",x"f5",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"ff",x"ff",x"ff",x"db",x"b7",x"92",x"6d",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"45",x"69",x"92",x"b6",x"d7",x"db",x"fb",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"db",x"b7",x"92",x"6e",x"49",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"24",x"24",x"49",x"49",x"6d",x"6d",x"6e",x"92",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"b6",x"ff",x"ff",x"ff",x"ff",x"ff",x"bb",x"71",x"04",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"29",x"49",x"49",x"6d",x"6d",x"8e",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"92",x"92",x"91",x"6d",x"49",x"48",x"24",x"00",x"00",x"00",x"00",x"45",x"92",x"db",x"db",x"db",x"db",x"fb",x"ff",x"ff",x"fb",x"fb",x"fb",x"db",x"db",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"db",x"fb",x"ff",x"ff",x"db",x"92",x"49",x"00",x"00",x"00",x"24",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"24",x"24",x"00",x"00",x"20",x"40",x"60",x"a4",x"c0",x"e0",x"e4",x"e0",x"e0",x"c0",x"c4",x"c9",x"f7",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"45",x"00",x"00",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"49",x"8e",x"b2",x"b7",x"db",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"db",x"b6",x"92",x"6e",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"6d",x"92",x"b6",x"db",x"db",x"fb",x"fb",x"fb",x"ff",x"ff",x"ff",x"fb",x"db",x"db",x"db",x"db",x"db",x"b2",x"6d",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"25",x"8e",x"ff",x"ff",x"ff",x"d6",x"ad",x"ac",x"cc",x"d0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f5",x"f1",x"f0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"f4",x"f5",x"f5",x"f5",x"fa",x"fa",x"fa",x"da",x"b6",x"6e",x"29",x"00",x"00",x"25",x"6d",x"92",x"d6",x"da",x"fb",x"fb",x"fa",x"fa",x"fa",x"f6",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fb",x"fb",x"db",x"b6",x"6e",x"49",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"48",x"49",x"69",x"6d",x"6e",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b7",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"6d",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"b6",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"df",x"96",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"24",x"49",x"49",x"69",x"6d",x"92",x"92",x"96",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"6d",x"6d",x"6d",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"b6",x"ff",x"ff",x"ff",x"fa",x"fa",x"fe",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"f9",x"f9",x"f5",x"f5",x"f6",x"f6",x"d6",x"b6",x"d6",x"ff",x"ff",x"ff",x"92",x"45",x"00",x"00",x"00",x"24",x"25",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"20",x"60",x"a4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"c9",x"f2",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"b6",x"24",x"00",x"20",x"24",x"48",x"49",x"28",x"28",x"49",x"29",x"25",x"25",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"49",x"8e",x"b6",x"db",x"fb",x"fb",x"fb",x"fa",x"fa",x"fa",x"fa",x"fa",x"f6",x"f6",x"f6",x"f6",x"f6",x"f6",x"fa",x"fa",x"fa",x"fa",x"fb",x"fb",x"db",x"b6",x"72",x"49",x"05",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"6e",x"92",x"b7",x"db",x"ff",x"ff",x"ff",x"fe",x"fa",x"fa",x"fa",x"f6",x"f6",x"f6",x"f6",x"f6",x"f6",x"f6",x"f6",x"fa",x"fb",x"ff",x"fb",x"db",x"bb",x"92",x"69",x"45",x"00",x"00",x"00",x"00",x"00",x"04",x"24",x"49",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"29",x"b7",x"ff",x"ff",x"fb",x"d6",x"ad",x"ac",x"ac",x"cc",x"cc",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f5",x"f9",x"fa",x"fa",x"fb",x"db",x"b6",x"6e",x"6e",x"92",x"d6",x"fb",x"fb",x"fa",x"fa",x"f6",x"f6",x"f1",x"f1",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f4",x"f4",x"f4",x"f5",x"f5",x"f5",x"f5",x"f9",x"fa",x"fa",x"ff",x"ff",x"fb",x"d7",x"b6",x"6e",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"44",x"49",x"6d",x"6e",x"6e",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"6d",x"6d",x"6d",x"49",x"6d",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"df",x"df",x"96",x"6d",x"49",x"49",x"49",x"29",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"45",x"49",x"69",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"92",x"71",x"6d",x"6d",x"69",x"45",x"24",x"00",x"00",x"00",x"00",x"49",x"db",x"ff",x"ff",x"fa",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f5",x"f5",x"f4",x"f4",x"f0",x"f0",x"f1",x"f1",x"8d",x"8d",x"b6",x"ff",x"ff",x"ff",x"6e",x"24",x"00",x"00",x"00",x"24",x"25",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"49",x"29",x"24",x"24",x"00",x"00",x"00",x"40",x"84",x"c4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e9",x"f2",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"8d",x"00",x"00",x"00",x"24",x"28",x"48",x"28",x"28",x"28",x"25",x"25",x"24",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"6d",x"b6",x"db",x"ff",x"ff",x"fe",x"fa",x"fa",x"f9",x"f9",x"f5",x"f5",x"f5",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f5",x"f5",x"f5",x"f6",x"fa",x"fa",x"fb",x"fb",x"db",x"b7",x"6e",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"6d",x"92",x"d7",x"df",x"ff",x"ff",x"fe",x"fe",x"fe",x"fe",x"f9",x"f9",x"f5",x"f0",x"f0",x"f1",x"f1",x"f1",x"f1",x"f1",x"f1",x"f5",x"f6",x"fa",x"fb",x"ff",x"ff",x"fb",x"d7",x"b2",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"6e",x"b7",x"ff",x"ff",x"ff",x"d6",x"b1",x"8c",x"88",x"ac",x"ac",x"d0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"f1",x"f5",x"f5",x"fa",x"fb",x"ff",x"fb",x"fb",x"fb",x"fb",x"f6",x"f6",x"f1",x"ed",x"ed",x"cc",x"cc",x"c8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f4",x"f4",x"f4",x"f5",x"d5",x"f5",x"f5",x"fa",x"fa",x"fb",x"ff",x"fb",x"b2",x"69",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"4d",x"6d",x"6d",x"6e",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"49",x"24",x"00",x"00",x"49",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"92",x"6d",x"6d",x"44",x"20",x"00",x"00",x"20",x"24",x"49",x"49",x"6d",x"6d",x"71",x"92",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"71",x"6d",x"69",x"49",x"24",x"00",x"00",x"00",x"00",x"25",x"6e",x"ff",x"ff",x"f9",x"f5",x"d5",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"d0",x"f0",x"f0",x"ec",x"ec",x"ec",x"cc",x"64",x"68",x"b6",x"ff",x"ff",x"db",x"49",x"00",x"00",x"00",x"00",x"24",x"45",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"29",x"24",x"24",x"00",x"00",x"00",x"20",x"60",x"a4",x"c4",x"e4",x"e0",x"e0",x"e0",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"c9",x"f2",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"8d",x"69",x"24",x"00",x"00",x"00",x"24",x"24",x"28",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"6e",x"b6",x"db",x"ff",x"ff",x"fe",x"fa",x"f9",x"f5",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f1",x"f1",x"d1",x"f6",x"fa",x"fb",x"ff",x"fb",x"b2",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"6d",x"b6",x"db",x"ff",x"ff",x"fe",x"fa",x"f9",x"f5",x"f5",x"f5",x"f4",x"f4",x"f4",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"cc",x"cc",x"ec",x"f1",x"f1",x"f5",x"f5",x"fa",x"fb",x"fb",x"d6",x"6d",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"6d",x"6d",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"04",x"00",x"00",x"00",x"00",x"00",x"49",x"92",x"ff",x"ff",x"ff",x"fb",x"d6",x"b1",x"8d",x"8c",x"88",x"88",x"a8",x"cc",x"cc",x"ec",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"d0",x"f1",x"f5",x"fa",x"fb",x"fa",x"f6",x"f1",x"cd",x"cc",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f5",x"f5",x"f5",x"f9",x"fa",x"fb",x"d7",x"92",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"28",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"24",x"00",x"00",x"49",x"b6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"d2",x"89",x"60",x"20",x"00",x"00",x"04",x"24",x"49",x"49",x"69",x"6d",x"92",x"96",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"6d",x"6d",x"49",x"45",x"24",x"00",x"00",x"00",x"00",x"49",x"b6",x"ff",x"fe",x"f9",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"ec",x"f0",x"f0",x"ec",x"ec",x"cc",x"a8",x"64",x"8d",x"da",x"ff",x"db",x"92",x"24",x"00",x"00",x"00",x"00",x"24",x"25",x"49",x"49",x"49",x"4d",x"6d",x"49",x"49",x"29",x"24",x"24",x"04",x"00",x"00",x"00",x"40",x"80",x"a4",x"e4",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c4",x"c9",x"f2",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"d2",x"89",x"44",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"6e",x"b7",x"ff",x"ff",x"ff",x"fe",x"f9",x"f9",x"f8",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"f0",x"f1",x"f1",x"f6",x"fb",x"ff",x"b6",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"92",x"db",x"ff",x"fe",x"fa",x"f9",x"f9",x"f9",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"d1",x"f6",x"fa",x"fb",x"d6",x"6d",x"24",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"24",x"04",x"00",x"00",x"00",x"00",x"00",x"49",x"92",x"db",x"ff",x"ff",x"ff",x"da",x"d6",x"b1",x"8d",x"88",x"88",x"88",x"a8",x"a8",x"a8",x"cc",x"cc",x"cc",x"cc",x"cc",x"cc",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"cc",x"cc",x"f0",x"f1",x"f5",x"f5",x"f1",x"cc",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f5",x"fb",x"fb",x"db",x"8e",x"25",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"24",x"00",x"00",x"24",x"6d",x"b6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f2",x"ee",x"c5",x"80",x"40",x"00",x"00",x"00",x"04",x"24",x"49",x"49",x"6d",x"71",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"49",x"49",x"25",x"20",x"00",x"00",x"00",x"04",x"92",x"db",x"ff",x"fa",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"ec",x"f0",x"ec",x"ec",x"ec",x"c8",x"84",x"88",x"b2",x"ff",x"ff",x"b7",x"49",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"4d",x"49",x"49",x"24",x"24",x"04",x"00",x"00",x"00",x"20",x"60",x"a0",x"c4",x"e4",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c4",x"c9",x"d2",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fa",x"d2",x"a9",x"85",x"64",x"20",x"00",x"00",x"00",x"00",x"04",x"24",x"24",x"24",x"25",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"8e",x"db",x"ff",x"ff",x"fe",x"fe",x"f9",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"f1",x"f6",x"fb",x"fb",x"b6",x"49",x"00",x"00",x"00",x"00",x"24",x"6e",x"b7",x"fb",x"ff",x"ff",x"fe",x"f9",x"f8",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"cc",x"d1",x"f5",x"fa",x"fb",x"d7",x"6d",x"04",x"00",x"00",x"00",x"24",x"24",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"72",x"db",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"b1",x"ad",x"8c",x"88",x"64",x"64",x"64",x"88",x"88",x"a8",x"a8",x"ac",x"cc",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"cc",x"cc",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"d0",x"d1",x"fa",x"ff",x"db",x"8e",x"25",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"92",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"ed",x"c9",x"c0",x"c0",x"c0",x"60",x"20",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"91",x"6d",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"49",x"b6",x"ff",x"fe",x"f9",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"a4",x"84",x"ad",x"fa",x"ff",x"ff",x"92",x"25",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"04",x"04",x"00",x"00",x"20",x"40",x"80",x"c4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"c9",x"f7",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"ce",x"a9",x"64",x"40",x"20",x"00",x"00",x"00",x"24",x"24",x"04",x"04",x"04",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"b2",x"db",x"ff",x"fe",x"f9",x"f9",x"d8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"c8",x"cd",x"f6",x"fb",x"fb",x"92",x"25",x"00",x"00",x"25",x"6e",x"db",x"ff",x"ff",x"fe",x"f9",x"f9",x"f8",x"f8",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"f0",x"ec",x"ec",x"ec",x"cc",x"cc",x"cc",x"d1",x"fa",x"ff",x"b6",x"49",x"00",x"00",x"00",x"00",x"24",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"44",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"05",x"49",x"72",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"da",x"d6",x"d6",x"b1",x"b1",x"8d",x"8d",x"88",x"88",x"88",x"88",x"88",x"ac",x"ac",x"ac",x"cc",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"e8",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c8",x"c8",x"c8",x"cc",x"ec",x"ec",x"f0",x"f0",x"f0",x"f0",x"f0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"ec",x"ec",x"ac",x"d1",x"fa",x"ff",x"db",x"6e",x"00",x"00",x"00",x"00",x"00",x"04",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"6d",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"ff",x"ff",x"ff",x"ff",x"fb",x"f2",x"e9",x"e5",x"e0",x"e0",x"e0",x"e0",x"a0",x"60",x"20",x"00",x"00",x"00",x"24",x"45",x"49",x"4d",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"00",x"00",x"00",x"04",x"92",x"db",x"ff",x"fa",x"f5",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"c8",x"84",x"64",x"d6",x"ff",x"ff",x"b7",x"4a",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"24",x"04",x"00",x"00",x"00",x"20",x"60",x"a4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"c0",x"a0",x"a9",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"ce",x"c9",x"c5",x"84",x"40",x"20",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"69",x"b6",x"ff",x"ff",x"fa",x"f9",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"c8",x"ad",x"f6",x"ff",x"db",x"4d",x"25",x"49",x"92",x"db",x"ff",x"fe",x"fa",x"f9",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"c8",x"cc",x"d6",x"ff",x"fb",x"92",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"6d",x"92",x"92",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"4d",x"49",x"44",x"48",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"6d",x"b6",x"b7",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"da",x"da",x"b6",x"b2",x"b2",x"91",x"8d",x"8c",x"8c",x"8c",x"ac",x"cc",x"d0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"e8",x"ec",x"ec",x"e8",x"c8",x"c4",x"a4",x"a4",x"a4",x"a8",x"a8",x"88",x"a8",x"c8",x"cc",x"ec",x"ec",x"f0",x"f0",x"f0",x"f0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"ec",x"ec",x"ec",x"cc",x"ac",x"d1",x"ff",x"ff",x"b7",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"b6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f2",x"e9",x"e5",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"40",x"20",x"00",x"00",x"24",x"24",x"49",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"49",x"49",x"44",x"24",x"00",x"00",x"00",x"25",x"d7",x"ff",x"fe",x"f9",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"cc",x"a8",x"64",x"89",x"db",x"ff",x"ff",x"92",x"25",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"24",x"24",x"04",x"00",x"00",x"20",x"40",x"84",x"c4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"c0",x"a4",x"a9",x"ad",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f2",x"cd",x"c9",x"a5",x"a0",x"60",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"69",x"b6",x"ff",x"ff",x"fe",x"d9",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"c8",x"a8",x"d2",x"fb",x"ff",x"92",x"6e",x"b7",x"db",x"ff",x"fe",x"f9",x"f8",x"f4",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f0",x"f0",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"c8",x"a8",x"b1",x"fb",x"ff",x"bb",x"25",x"00",x"00",x"00",x"24",x"24",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"44",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"6e",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"db",x"d6",x"d6",x"b1",x"b1",x"b0",x"cc",x"cc",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"c8",x"a8",x"84",x"60",x"60",x"40",x"44",x"64",x"68",x"88",x"a8",x"a8",x"a8",x"cc",x"ec",x"ec",x"f0",x"f0",x"f0",x"f0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ac",x"ac",x"fa",x"ff",x"db",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"b6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d2",x"c5",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"a4",x"80",x"40",x"00",x"00",x"00",x"24",x"24",x"44",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"48",x"24",x"00",x"00",x"00",x"00",x"6d",x"fb",x"ff",x"fa",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"cc",x"84",x"88",x"b2",x"ff",x"ff",x"db",x"49",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"48",x"44",x"24",x"24",x"00",x"00",x"00",x"20",x"80",x"c4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"c0",x"a0",x"a9",x"b1",x"d6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f2",x"c9",x"a5",x"a5",x"80",x"60",x"40",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"d7",x"ff",x"ff",x"fa",x"f9",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"ec",x"cc",x"a8",x"ad",x"d6",x"ff",x"db",x"db",x"fb",x"fb",x"fa",x"f9",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"c8",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"ec",x"ec",x"a8",x"ad",x"fb",x"ff",x"db",x"49",x"00",x"00",x"00",x"24",x"24",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"44",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"49",x"6e",x"92",x"b7",x"db",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fa",x"d6",x"d1",x"b0",x"d0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"c8",x"84",x"60",x"64",x"68",x"8d",x"91",x"b2",x"b2",x"b6",x"d6",x"d1",x"cd",x"cd",x"cd",x"ec",x"ec",x"f0",x"f0",x"f0",x"f0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"a8",x"a8",x"f6",x"ff",x"db",x"6e",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"b6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"d7",x"ad",x"a5",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"60",x"20",x"00",x"00",x"00",x"04",x"24",x"49",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"6d",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"49",x"92",x"ff",x"ff",x"f9",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"cc",x"a8",x"68",x"8d",x"da",x"ff",x"df",x"97",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"20",x"60",x"a0",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a5",x"ad",x"b6",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d2",x"a9",x"a5",x"84",x"60",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"b2",x"fb",x"ff",x"fa",x"f9",x"f4",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"c8",x"a4",x"80",x"80",x"a4",x"c4",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"ec",x"c8",x"88",x"8d",x"d6",x"ff",x"ff",x"ff",x"fb",x"fa",x"f9",x"f4",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"e8",x"c8",x"a8",x"84",x"80",x"a4",x"c4",x"c8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"84",x"88",x"d6",x"ff",x"ff",x"6e",x"24",x"00",x"00",x"20",x"24",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"49",x"6e",x"92",x"92",x"96",x"b7",x"db",x"db",x"db",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"da",x"d5",x"d0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"c8",x"a4",x"64",x"64",x"69",x"92",x"da",x"df",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"d6",x"d1",x"d1",x"f0",x"f0",x"f0",x"f0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"a8",x"a8",x"d6",x"fb",x"ff",x"92",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"ae",x"a5",x"c4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"40",x"20",x"00",x"00",x"00",x"24",x"45",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"df",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"28",x"24",x"00",x"00",x"00",x"00",x"6e",x"db",x"ff",x"fa",x"f5",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"c8",x"88",x"88",x"b2",x"ff",x"ff",x"db",x"6e",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"28",x"24",x"24",x"20",x"00",x"00",x"00",x"20",x"64",x"c4",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"c1",x"c5",x"a9",x"b2",x"bb",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d2",x"a9",x"84",x"60",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"92",x"fb",x"ff",x"fa",x"f9",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"c8",x"a4",x"84",x"64",x"84",x"88",x"a8",x"c8",x"e8",x"e8",x"e8",x"ec",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"a8",x"84",x"ad",x"da",x"ff",x"ff",x"fe",x"fa",x"f9",x"f4",x"f4",x"f4",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"a8",x"84",x"64",x"84",x"84",x"a8",x"c8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"c8",x"84",x"68",x"d6",x"ff",x"df",x"72",x"24",x"00",x"00",x"00",x"24",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"6e",x"72",x"97",x"db",x"ff",x"ff",x"ff",x"ff",x"da",x"f1",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"c8",x"84",x"60",x"64",x"b1",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"d5",x"d0",x"f0",x"f0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"a4",x"84",x"d6",x"ff",x"ff",x"92",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"92",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"b6",x"ad",x"a5",x"c4",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"c0",x"60",x"20",x"00",x"00",x"00",x"24",x"44",x"49",x"49",x"6d",x"92",x"92",x"92",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"24",x"b6",x"ff",x"ff",x"f6",x"f0",x"f0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"a8",x"88",x"8d",x"b6",x"ff",x"ff",x"b6",x"45",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"28",x"24",x"24",x"20",x"00",x"00",x"00",x"40",x"84",x"e5",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"c4",x"c1",x"a9",x"ae",x"b6",x"bb",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"d6",x"89",x"40",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"20",x"20",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"92",x"db",x"ff",x"fa",x"f9",x"f8",x"f8",x"f8",x"f4",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"ec",x"ec",x"e8",x"e8",x"e8",x"a4",x"84",x"64",x"8d",x"b2",x"d6",x"d2",x"cd",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c8",x"a4",x"64",x"d1",x"ff",x"ff",x"ff",x"fa",x"f9",x"f8",x"f8",x"f4",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"e8",x"e8",x"c8",x"a8",x"84",x"88",x"d2",x"d6",x"d2",x"d1",x"cc",x"cc",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"e8",x"a4",x"84",x"8d",x"fb",x"ff",x"df",x"4d",x"24",x"00",x"00",x"20",x"24",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"6d",x"4d",x"49",x"24",x"24",x"24",x"44",x"44",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"69",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"25",x"49",x"6e",x"b7",x"db",x"ff",x"ff",x"fa",x"f5",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"e8",x"a4",x"44",x"68",x"b2",x"db",x"ff",x"ff",x"ff",x"db",x"bb",x"b7",x"b7",x"b7",x"db",x"ff",x"ff",x"fa",x"f5",x"d0",x"f0",x"f0",x"f0",x"f0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"84",x"64",x"d6",x"ff",x"ff",x"92",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"49",x"69",x"6d",x"6e",x"6e",x"8e",x"8e",x"6e",x"6d",x"6d",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"b6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"df",x"bb",x"92",x"89",x"a5",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"c0",x"a0",x"40",x"00",x"00",x"00",x"20",x"24",x"29",x"49",x"69",x"6d",x"92",x"92",x"b6",x"b6",x"ba",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"4d",x"db",x"ff",x"fa",x"f5",x"f0",x"f0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"cc",x"84",x"64",x"b6",x"df",x"ff",x"db",x"6e",x"00",x"00",x"00",x"00",x"04",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"44",x"44",x"24",x"00",x"00",x"00",x"00",x"20",x"84",x"c4",x"e4",x"e0",x"e0",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"c0",x"a4",x"a9",x"ae",x"b6",x"bb",x"bf",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"d6",x"49",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"4a",x"db",x"ff",x"fe",x"f9",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"ec",x"ec",x"e8",x"ec",x"e8",x"c8",x"80",x"64",x"b2",x"d7",x"ff",x"ff",x"fa",x"f1",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"a4",x"84",x"88",x"d6",x"ff",x"ff",x"fa",x"f9",x"f9",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"e8",x"e8",x"c8",x"a4",x"64",x"8d",x"d6",x"ff",x"ff",x"fa",x"f1",x"ec",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"e8",x"ec",x"c8",x"84",x"88",x"b2",x"ff",x"ff",x"b7",x"45",x"00",x"00",x"00",x"24",x"44",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"4d",x"49",x"28",x"24",x"04",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"44",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"92",x"db",x"ff",x"fe",x"f5",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f4",x"f4",x"f0",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"e8",x"c4",x"84",x"48",x"92",x"db",x"ff",x"ff",x"db",x"b7",x"92",x"6d",x"49",x"49",x"6e",x"92",x"b7",x"ff",x"fa",x"f5",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"c8",x"64",x"64",x"fb",x"ff",x"ff",x"72",x"25",x"00",x"00",x"00",x"00",x"20",x"25",x"49",x"92",x"b6",x"d7",x"db",x"db",x"fb",x"fb",x"fb",x"fb",x"db",x"d6",x"b2",x"6e",x"45",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"da",x"ff",x"ff",x"ff",x"ff",x"df",x"df",x"df",x"df",x"df",x"ff",x"ff",x"ff",x"ff",x"df",x"df",x"bf",x"96",x"92",x"89",x"a5",x"c0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"c4",x"80",x"20",x"00",x"00",x"00",x"20",x"24",x"29",x"49",x"6d",x"8d",x"92",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"91",x"6d",x"49",x"49",x"24",x"20",x"00",x"00",x"00",x"24",x"92",x"ff",x"ff",x"f6",x"f1",x"f0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"a8",x"64",x"68",x"da",x"ff",x"ff",x"92",x"25",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"29",x"44",x"44",x"24",x"00",x"00",x"00",x"00",x"40",x"a4",x"e4",x"e0",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c4",x"c4",x"a5",x"8e",x"96",x"9b",x"9f",x"bf",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"d7",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"92",x"ff",x"ff",x"f9",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"ec",x"ec",x"ec",x"ec",x"e8",x"ec",x"e8",x"c4",x"60",x"69",x"db",x"ff",x"ff",x"ff",x"fa",x"f1",x"e8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"c8",x"a4",x"84",x"ad",x"fb",x"ff",x"ff",x"f9",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"a8",x"84",x"68",x"b6",x"ff",x"ff",x"ff",x"ff",x"f1",x"ec",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"a8",x"64",x"8d",x"b6",x"ff",x"ff",x"b2",x"24",x"00",x"00",x"00",x"24",x"49",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"6d",x"49",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"24",x"24",x"24",x"24",x"28",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6a",x"b7",x"ff",x"fa",x"f5",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f4",x"f4",x"f0",x"f4",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"c8",x"80",x"84",x"b2",x"db",x"ff",x"ff",x"db",x"8e",x"49",x"24",x"00",x"00",x"00",x"00",x"25",x"92",x"fb",x"fb",x"f9",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"a8",x"88",x"8d",x"fb",x"ff",x"df",x"29",x"00",x"00",x"00",x"25",x"49",x"b2",x"d7",x"db",x"fb",x"ff",x"ff",x"ff",x"fe",x"fe",x"fe",x"fe",x"fe",x"fa",x"fa",x"fb",x"fb",x"d7",x"92",x"49",x"24",x"00",x"00",x"00",x"00",x"20",x"6d",x"db",x"ff",x"df",x"df",x"bf",x"bf",x"9f",x"9b",x"96",x"b6",x"d7",x"fb",x"ff",x"ff",x"ff",x"df",x"bf",x"9b",x"97",x"92",x"a9",x"c4",x"e0",x"e0",x"e0",x"e4",x"e0",x"e0",x"e0",x"e0",x"a0",x"60",x"20",x"00",x"00",x"00",x"04",x"24",x"49",x"69",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"4d",x"db",x"ff",x"fa",x"f5",x"f0",x"f0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"c8",x"84",x"84",x"8d",x"db",x"ff",x"df",x"6d",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"44",x"24",x"00",x"00",x"00",x"00",x"20",x"80",x"a0",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c4",x"c5",x"a9",x"92",x"77",x"9b",x"bf",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"df",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"d6",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"6d",x"d7",x"ff",x"fe",x"f9",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"c8",x"a4",x"84",x"ad",x"fb",x"ff",x"ff",x"fe",x"f5",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c8",x"84",x"88",x"d6",x"ff",x"ff",x"fe",x"f9",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"a4",x"84",x"ad",x"da",x"ff",x"ff",x"ff",x"fa",x"ed",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c8",x"a8",x"84",x"b1",x"db",x"ff",x"db",x"92",x"20",x"00",x"00",x"00",x"24",x"49",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"00",x"00",x"00",x"49",x"4d",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"24",x"24",x"24",x"24",x"24",x"45",x"28",x"28",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6a",x"d7",x"ff",x"fa",x"f5",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"c8",x"a8",x"84",x"84",x"da",x"ff",x"ff",x"db",x"8e",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"72",x"ff",x"ff",x"f5",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"c8",x"84",x"88",x"b2",x"ff",x"ff",x"b7",x"01",x"00",x"25",x"69",x"92",x"d7",x"db",x"fa",x"fe",x"fe",x"fe",x"fa",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fa",x"fa",x"fa",x"fb",x"fb",x"b7",x"6e",x"20",x"00",x"00",x"00",x"24",x"92",x"ff",x"ff",x"bf",x"9f",x"7f",x"7f",x"7b",x"7b",x"77",x"72",x"92",x"d2",x"f6",x"fb",x"ff",x"ff",x"df",x"9b",x"7b",x"77",x"92",x"a9",x"c0",x"e0",x"e0",x"e4",x"e0",x"e0",x"e0",x"e0",x"c4",x"a0",x"40",x"00",x"00",x"00",x"00",x"24",x"29",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"b7",x"b6",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"25",x"92",x"ff",x"ff",x"fa",x"f5",x"f0",x"f0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"c8",x"60",x"89",x"d6",x"ff",x"ff",x"bb",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"60",x"a4",x"c0",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e0",x"e0",x"e0",x"c0",x"c5",x"c9",x"ae",x"77",x"7b",x"9b",x"bf",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"d6",x"b6",x"9b",x"9b",x"bf",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"d6",x"69",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"b2",x"ff",x"ff",x"fa",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"a4",x"80",x"ad",x"d6",x"ff",x"ff",x"ff",x"fa",x"f1",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"a4",x"84",x"ad",x"fa",x"ff",x"ff",x"fa",x"f5",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"c8",x"80",x"84",x"d6",x"ff",x"ff",x"ff",x"fb",x"f6",x"cc",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"a8",x"84",x"88",x"d6",x"ff",x"ff",x"b7",x"49",x"00",x"00",x"00",x"04",x"24",x"49",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"24",x"00",x"00",x"00",x"29",x"96",x"bb",x"96",x"29",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"28",x"28",x"28",x"28",x"29",x"49",x"49",x"49",x"49",x"44",x"44",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"8e",x"db",x"ff",x"fa",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"c8",x"84",x"84",x"8d",x"fb",x"ff",x"ff",x"8e",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"29",x"97",x"ff",x"fa",x"f5",x"f0",x"f0",x"f0",x"f0",x"f0",x"f4",x"f0",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"a4",x"44",x"8d",x"fa",x"ff",x"ff",x"93",x"25",x"25",x"6e",x"b6",x"fb",x"ff",x"fe",x"f9",x"f9",x"f9",x"f9",x"f4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f4",x"f0",x"d0",x"f5",x"f6",x"fb",x"fb",x"d7",x"49",x"00",x"00",x"00",x"49",x"bb",x"df",x"bf",x"9f",x"7f",x"5f",x"5b",x"5b",x"7b",x"7b",x"77",x"72",x"8d",x"ad",x"d2",x"fb",x"ff",x"df",x"7b",x"5b",x"7b",x"97",x"ae",x"a4",x"c0",x"e0",x"e4",x"e0",x"e0",x"e0",x"e0",x"e4",x"c4",x"80",x"20",x"00",x"00",x"00",x"04",x"24",x"49",x"49",x"6d",x"6d",x"92",x"92",x"b2",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"6e",x"db",x"ff",x"fa",x"f5",x"f4",x"f0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"c8",x"a4",x"64",x"b1",x"fb",x"ff",x"db",x"72",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"04",x"00",x"00",x"00",x"40",x"80",x"c4",x"e0",x"e0",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"c0",x"c4",x"a9",x"ae",x"92",x"7b",x"7b",x"9f",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"f6",x"f2",x"ae",x"8e",x"72",x"76",x"7b",x"9b",x"df",x"ff",x"ff",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"6d",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"8e",x"db",x"ff",x"fa",x"f5",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"c4",x"a4",x"64",x"b2",x"ff",x"ff",x"ff",x"ff",x"f6",x"ec",x"c4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"84",x"88",x"b2",x"ff",x"ff",x"fe",x"f9",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"a4",x"60",x"88",x"db",x"ff",x"ff",x"ff",x"fa",x"f1",x"c8",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"84",x"84",x"ad",x"fb",x"ff",x"df",x"6e",x"24",x"00",x"00",x"00",x"24",x"24",x"49",x"4d",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"44",x"20",x"00",x"00",x"4d",x"bb",x"df",x"df",x"9b",x"9b",x"77",x"56",x"2d",x"09",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"44",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"d7",x"ff",x"fa",x"f5",x"f0",x"ec",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"c8",x"64",x"88",x"b6",x"ff",x"ff",x"b6",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"72",x"df",x"ff",x"fa",x"f1",x"ec",x"f0",x"f0",x"f0",x"f0",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"c8",x"a4",x"68",x"b6",x"ff",x"ff",x"b7",x"92",x"92",x"b6",x"ff",x"ff",x"fa",x"fa",x"f9",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"ec",x"ec",x"cc",x"d0",x"d1",x"fb",x"fb",x"b3",x"49",x"00",x"00",x"4d",x"bf",x"bf",x"9b",x"5b",x"5b",x"5f",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"8e",x"89",x"84",x"cd",x"f6",x"fb",x"9b",x"7b",x"5b",x"77",x"92",x"8d",x"a4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c4",x"c4",x"a0",x"60",x"20",x"00",x"00",x"00",x"24",x"28",x"49",x"4d",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"25",x"92",x"fb",x"ff",x"fa",x"f4",x"f0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"a8",x"84",x"88",x"d6",x"ff",x"ff",x"97",x"29",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"04",x"00",x"00",x"00",x"20",x"60",x"a4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"c0",x"a5",x"8d",x"92",x"97",x"5b",x"7f",x"bf",x"df",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"d2",x"a9",x"a9",x"a9",x"89",x"92",x"7b",x"7f",x"5b",x"7b",x"97",x"bb",x"bf",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"b2",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"b7",x"ff",x"ff",x"f9",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"a0",x"80",x"89",x"da",x"ff",x"ff",x"ff",x"fa",x"f1",x"e8",x"e4",x"e4",x"e4",x"e8",x"e8",x"e8",x"e4",x"e8",x"a4",x"64",x"8d",x"da",x"ff",x"fe",x"fa",x"f5",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"c8",x"84",x"84",x"ad",x"fb",x"ff",x"ff",x"fb",x"f6",x"ed",x"c8",x"c4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c8",x"64",x"68",x"d6",x"ff",x"ff",x"bb",x"29",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"6d",x"6d",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"04",x"92",x"ff",x"ff",x"bf",x"9b",x"9b",x"7b",x"7b",x"57",x"32",x"32",x"29",x"05",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"28",x"29",x"28",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"92",x"fb",x"ff",x"fa",x"f5",x"f0",x"ec",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"c8",x"88",x"64",x"b1",x"da",x"ff",x"db",x"6e",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"b7",x"ff",x"ff",x"f5",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"c8",x"a4",x"84",x"8d",x"da",x"ff",x"df",x"b7",x"b6",x"db",x"ff",x"ff",x"fa",x"f9",x"f5",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"ec",x"ec",x"f0",x"cc",x"ac",x"ac",x"d6",x"fb",x"fb",x"92",x"05",x"00",x"29",x"9b",x"9b",x"7b",x"5b",x"5b",x"5b",x"5f",x"3f",x"5f",x"5b",x"5f",x"7b",x"96",x"8d",x"65",x"84",x"c9",x"d2",x"b6",x"97",x"7b",x"7b",x"77",x"92",x"a9",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c4",x"e4",x"c4",x"a0",x"60",x"20",x"00",x"00",x"24",x"24",x"29",x"49",x"4d",x"6d",x"8d",x"92",x"92",x"92",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"d7",x"fb",x"fa",x"f5",x"f0",x"f0",x"f4",x"f4",x"f0",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"e8",x"ec",x"ec",x"84",x"84",x"ad",x"fb",x"ff",x"db",x"6e",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"40",x"84",x"c4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e0",x"e0",x"c0",x"a4",x"a9",x"92",x"7b",x"7b",x"5b",x"9f",x"df",x"ff",x"ff",x"fb",x"fa",x"f6",x"d1",x"ed",x"c9",x"a0",x"a4",x"89",x"8e",x"76",x"7b",x"5f",x"5f",x"5b",x"5b",x"7b",x"9b",x"9f",x"bf",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"da",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"db",x"ff",x"fe",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"c8",x"80",x"84",x"b1",x"fb",x"ff",x"ff",x"ff",x"f6",x"ed",x"e8",x"e4",x"e4",x"e4",x"e4",x"e8",x"e8",x"e4",x"c4",x"80",x"84",x"b6",x"ff",x"ff",x"fe",x"f9",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"a4",x"84",x"ad",x"d6",x"ff",x"ff",x"ff",x"fa",x"f1",x"e8",x"e8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"a4",x"64",x"8d",x"db",x"ff",x"df",x"72",x"25",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"6d",x"6d",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"4d",x"b6",x"ff",x"df",x"bf",x"7b",x"5b",x"5b",x"5f",x"7f",x"7f",x"5b",x"57",x"4e",x"29",x"05",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"29",x"b7",x"ff",x"ff",x"f5",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"e8",x"e8",x"e8",x"c8",x"84",x"64",x"89",x"b6",x"ff",x"ff",x"b7",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"db",x"ff",x"fa",x"d1",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"c8",x"84",x"88",x"b6",x"db",x"ff",x"ff",x"db",x"fb",x"ff",x"fa",x"f9",x"f5",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"f0",x"ec",x"cc",x"88",x"b1",x"fb",x"ff",x"b7",x"25",x"00",x"05",x"2e",x"77",x"7b",x"7b",x"5b",x"5b",x"3b",x"3f",x"3f",x"5f",x"5f",x"7f",x"7b",x"96",x"8d",x"84",x"a4",x"a5",x"ae",x"92",x"97",x"77",x"7b",x"7b",x"92",x"a9",x"c5",x"e0",x"e0",x"e0",x"e0",x"c0",x"e4",x"c4",x"c4",x"80",x"40",x"00",x"00",x"00",x"04",x"28",x"49",x"49",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"25",x"92",x"fb",x"fb",x"f6",x"f5",x"f0",x"f0",x"f0",x"f4",x"f0",x"f0",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"e8",x"e8",x"cc",x"84",x"64",x"d6",x"ff",x"ff",x"b7",x"29",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"20",x"60",x"a4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e0",x"e0",x"c0",x"c4",x"a9",x"8e",x"76",x"7b",x"5f",x"7b",x"bf",x"ff",x"fb",x"f7",x"f2",x"ed",x"c9",x"c4",x"c4",x"c0",x"c0",x"a5",x"8e",x"96",x"7b",x"5f",x"5f",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"9f",x"bf",x"df",x"df",x"ff",x"ff",x"ff",x"db",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"b6",x"ff",x"ff",x"f9",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"c4",x"80",x"88",x"d6",x"ff",x"ff",x"ff",x"fa",x"f1",x"e8",x"e4",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"80",x"80",x"89",x"da",x"ff",x"fe",x"fa",x"f5",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"c4",x"84",x"84",x"d2",x"fb",x"ff",x"ff",x"ff",x"f6",x"ed",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"84",x"68",x"b2",x"ff",x"ff",x"db",x"49",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"24",x"ba",x"ff",x"ff",x"df",x"bf",x"9f",x"7b",x"5b",x"5f",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"77",x"52",x"2d",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"04",x"6e",x"fb",x"ff",x"fa",x"d1",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"c8",x"84",x"64",x"b2",x"fb",x"ff",x"db",x"6e",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"b6",x"ff",x"ff",x"f5",x"d0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"c8",x"a4",x"84",x"8d",x"db",x"ff",x"ff",x"db",x"ff",x"ff",x"fa",x"f5",x"f4",x"f0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"e8",x"ec",x"ec",x"cc",x"88",x"ad",x"fa",x"ff",x"b7",x"49",x"01",x"00",x"00",x"4e",x"77",x"9f",x"7f",x"5b",x"3b",x"3b",x"3f",x"5f",x"5b",x"5b",x"5b",x"7b",x"b6",x"ad",x"a9",x"a4",x"85",x"89",x"92",x"97",x"7b",x"7b",x"97",x"92",x"85",x"c0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"c4",x"a0",x"60",x"20",x"00",x"00",x"00",x"24",x"28",x"49",x"69",x"6d",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"db",x"ff",x"fa",x"f5",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"e8",x"c8",x"a8",x"84",x"8d",x"db",x"ff",x"df",x"6e",x"05",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"20",x"40",x"80",x"a4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c4",x"a5",x"8e",x"92",x"7b",x"5f",x"7f",x"9f",x"ba",x"d6",x"ee",x"e9",x"c4",x"c0",x"c0",x"c0",x"c0",x"c4",x"c5",x"ae",x"97",x"7b",x"5f",x"3f",x"3b",x"3b",x"3b",x"3f",x"3f",x"5f",x"7b",x"7b",x"9b",x"bf",x"bf",x"df",x"ff",x"ff",x"ff",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"db",x"ff",x"fa",x"f5",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"c8",x"a4",x"84",x"ad",x"ff",x"ff",x"ff",x"fb",x"f6",x"ed",x"c4",x"e4",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"c4",x"60",x"64",x"b2",x"ff",x"ff",x"fe",x"f5",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"a4",x"84",x"89",x"db",x"ff",x"ff",x"ff",x"fa",x"f1",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"a4",x"60",x"8d",x"db",x"ff",x"ff",x"92",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"24",x"24",x"24",x"00",x"00",x"24",x"6d",x"ff",x"ff",x"ff",x"ff",x"df",x"9f",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5f",x"7f",x"7f",x"7f",x"7b",x"56",x"52",x"2d",x"29",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"b6",x"ff",x"ff",x"f6",x"d0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"a8",x"64",x"69",x"db",x"ff",x"ff",x"b7",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"db",x"ff",x"fa",x"f5",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"c8",x"84",x"88",x"b1",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"f5",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"c8",x"a8",x"64",x"8d",x"da",x"ff",x"b7",x"49",x"01",x"00",x"00",x"04",x"4d",x"76",x"7b",x"5f",x"3b",x"3b",x"3b",x"5f",x"5b",x"5b",x"5b",x"7b",x"97",x"92",x"ae",x"a9",x"a4",x"85",x"ae",x"92",x"77",x"7b",x"7b",x"96",x"6d",x"a5",x"c0",x"e0",x"e0",x"e0",x"e0",x"c4",x"c4",x"a0",x"60",x"40",x"20",x"00",x"00",x"04",x"24",x"49",x"49",x"6d",x"6d",x"72",x"72",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"25",x"24",x"00",x"00",x"00",x"00",x"24",x"8e",x"ff",x"ff",x"fa",x"f5",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"c8",x"84",x"88",x"b2",x"ff",x"ff",x"db",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"20",x"60",x"80",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c4",x"a5",x"8d",x"92",x"77",x"7b",x"7b",x"7b",x"b6",x"b1",x"a9",x"c5",x"e0",x"c0",x"e0",x"e0",x"e4",x"c5",x"a9",x"ae",x"b7",x"9b",x"7f",x"5f",x"3b",x"3b",x"5b",x"5b",x"3f",x"3f",x"3b",x"5b",x"7b",x"7b",x"7f",x"9f",x"bf",x"df",x"ff",x"ff",x"6d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"92",x"ff",x"fa",x"f9",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"c8",x"a4",x"84",x"89",x"d2",x"ff",x"ff",x"ff",x"f6",x"f1",x"e8",x"e4",x"e4",x"e4",x"e4",x"e8",x"e8",x"e8",x"e4",x"a4",x"60",x"89",x"da",x"ff",x"ff",x"fa",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"c8",x"80",x"64",x"b2",x"fb",x"ff",x"ff",x"fb",x"f6",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"84",x"64",x"b6",x"ff",x"ff",x"db",x"6e",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"6d",x"6d",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"6d",x"da",x"ff",x"ff",x"ff",x"ff",x"df",x"bf",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5f",x"5f",x"5f",x"7f",x"7b",x"7b",x"77",x"2e",x"05",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"db",x"ff",x"fa",x"f1",x"cc",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"c8",x"a4",x"88",x"ad",x"ff",x"ff",x"fb",x"8e",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"92",x"ff",x"fe",x"f5",x"f1",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"a8",x"84",x"8d",x"d6",x"ff",x"ff",x"ff",x"ff",x"ff",x"fa",x"f1",x"f0",x"f0",x"f0",x"f0",x"ec",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"c8",x"84",x"64",x"ad",x"da",x"ff",x"b6",x"49",x"00",x"00",x"00",x"00",x"04",x"2d",x"56",x"7b",x"5b",x"5b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"77",x"92",x"ae",x"a9",x"a4",x"a9",x"8e",x"96",x"77",x"7b",x"7b",x"72",x"89",x"a5",x"e0",x"e0",x"e0",x"e0",x"c0",x"c4",x"c0",x"80",x"60",x"20",x"00",x"00",x"04",x"24",x"48",x"49",x"69",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"69",x"b6",x"ff",x"fa",x"f5",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"a8",x"64",x"8d",x"da",x"ff",x"ff",x"96",x"00",x"00",x"00",x"00",x"00",x"04",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"40",x"60",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"c0",x"c5",x"ad",x"92",x"77",x"7b",x"7b",x"77",x"72",x"a9",x"a4",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"c5",x"a9",x"8e",x"96",x"7b",x"7b",x"5b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5f",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"9f",x"bf",x"df",x"df",x"92",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"db",x"ff",x"fa",x"f5",x"f4",x"f4",x"f0",x"f0",x"f4",x"f4",x"f4",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"c4",x"84",x"64",x"b1",x"db",x"ff",x"ff",x"fa",x"f6",x"ed",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e8",x"c4",x"84",x"88",x"b2",x"ff",x"ff",x"fa",x"f5",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"c8",x"a4",x"64",x"89",x"d6",x"ff",x"ff",x"ff",x"fa",x"f1",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"a0",x"64",x"6d",x"db",x"ff",x"ff",x"92",x"25",x"00",x"00",x"00",x"00",x"04",x"24",x"44",x"49",x"49",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"28",x"b6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"bf",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"56",x"52",x"2e",x"29",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"b6",x"ff",x"fb",x"f6",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"c8",x"64",x"89",x"d6",x"ff",x"ff",x"d7",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6e",x"db",x"ff",x"fa",x"f1",x"d0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f4",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"a4",x"64",x"b1",x"db",x"ff",x"ff",x"ff",x"ff",x"fa",x"f5",x"d0",x"ec",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"a4",x"60",x"89",x"d6",x"ff",x"ff",x"b6",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"29",x"52",x"7b",x"7f",x"5f",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"97",x"b2",x"a9",x"a4",x"a4",x"89",x"92",x"77",x"7b",x"7b",x"77",x"92",x"89",x"c4",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"60",x"20",x"00",x"00",x"04",x"24",x"24",x"45",x"49",x"49",x"4d",x"4d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"92",x"ff",x"ff",x"fa",x"d4",x"d0",x"f0",x"f0",x"f0",x"f0",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"a8",x"68",x"b2",x"ff",x"ff",x"bb",x"6d",x"00",x"00",x"00",x"00",x"00",x"04",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"20",x"40",x"80",x"a4",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e4",x"e0",x"e0",x"c4",x"a9",x"8e",x"77",x"7b",x"7b",x"77",x"76",x"8e",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c4",x"c5",x"ae",x"96",x"7b",x"5f",x"5f",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3f",x"5b",x"5b",x"7b",x"9b",x"bf",x"ff",x"bb",x"6d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"92",x"ff",x"ff",x"f9",x"f4",x"f4",x"f0",x"f0",x"f0",x"f4",x"f4",x"f4",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"a4",x"64",x"64",x"d6",x"ff",x"ff",x"ff",x"fa",x"f1",x"e8",x"e4",x"e4",x"e4",x"e8",x"e4",x"e4",x"e4",x"e8",x"a4",x"60",x"8d",x"da",x"ff",x"ff",x"fa",x"f5",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"c8",x"a4",x"84",x"8d",x"db",x"ff",x"ff",x"ff",x"f6",x"cc",x"c8",x"e8",x"e8",x"e4",x"e8",x"c8",x"e8",x"e8",x"c4",x"80",x"84",x"b6",x"ff",x"ff",x"db",x"49",x"00",x"00",x"00",x"00",x"04",x"04",x"24",x"49",x"49",x"49",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"92",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"9b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7f",x"7f",x"7b",x"77",x"52",x"2e",x"29",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"db",x"ff",x"fa",x"f1",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"a4",x"64",x"ad",x"fb",x"ff",x"ff",x"92",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"21",x"b2",x"ff",x"ff",x"f5",x"f0",x"ec",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"c4",x"84",x"88",x"d6",x"ff",x"ff",x"ff",x"ff",x"ff",x"f6",x"d1",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"c8",x"a4",x"60",x"64",x"ae",x"db",x"ff",x"df",x"72",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"29",x"76",x"7b",x"7f",x"5b",x"3b",x"3b",x"5b",x"5b",x"5f",x"5b",x"7b",x"97",x"b2",x"a9",x"a5",x"89",x"89",x"92",x"77",x"77",x"7b",x"76",x"8d",x"a9",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"80",x"60",x"20",x"00",x"00",x"04",x"24",x"44",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"d7",x"ff",x"fa",x"f5",x"d0",x"cc",x"f0",x"f0",x"f0",x"f0",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"a4",x"84",x"8d",x"da",x"ff",x"ff",x"92",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"20",x"40",x"80",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e4",x"e0",x"c0",x"a5",x"8d",x"76",x"7b",x"7b",x"7b",x"92",x"8e",x"a9",x"c0",x"e0",x"e0",x"e0",x"e0",x"c4",x"c4",x"a9",x"ad",x"96",x"7b",x"5f",x"5f",x"3f",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"5b",x"7b",x"9f",x"df",x"bb",x"6d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"db",x"ff",x"ff",x"f5",x"f4",x"f4",x"f0",x"f0",x"f0",x"f4",x"f4",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"a0",x"64",x"89",x"db",x"ff",x"ff",x"ff",x"f6",x"ed",x"e4",x"e4",x"e4",x"e4",x"e8",x"e4",x"e4",x"e4",x"e4",x"a0",x"60",x"b2",x"df",x"ff",x"ff",x"f5",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"80",x"89",x"b6",x"ff",x"ff",x"ff",x"fa",x"f1",x"c8",x"c4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"80",x"8d",x"db",x"ff",x"ff",x"b6",x"25",x"00",x"00",x"00",x"00",x"04",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"71",x"92",x"92",x"92",x"8d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"29",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"bf",x"7b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5f",x"5f",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5f",x"7f",x"7f",x"7b",x"57",x"52",x"2d",x"05",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"92",x"ff",x"fe",x"f5",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"a4",x"84",x"88",x"d6",x"ff",x"ff",x"b7",x"4e",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"db",x"ff",x"fa",x"f1",x"ec",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"c8",x"80",x"84",x"b2",x"fb",x"ff",x"df",x"ff",x"ff",x"ff",x"d5",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"e8",x"c8",x"a8",x"40",x"44",x"8d",x"bb",x"df",x"df",x"97",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"29",x"52",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5f",x"3b",x"5b",x"7b",x"97",x"92",x"8d",x"85",x"a4",x"c9",x"92",x"77",x"57",x"57",x"76",x"8e",x"a5",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"80",x"60",x"20",x"00",x"00",x"00",x"24",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"25",x"24",x"00",x"00",x"00",x"00",x"04",x"6e",x"db",x"ff",x"fa",x"f5",x"d0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"c8",x"84",x"84",x"b6",x"ff",x"ff",x"db",x"6d",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"48",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"00",x"00",x"20",x"40",x"60",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"e0",x"e0",x"c0",x"c0",x"a4",x"89",x"72",x"5b",x"7f",x"7b",x"93",x"ae",x"a9",x"a4",x"c0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a9",x"8d",x"96",x"7b",x"7b",x"7f",x"3b",x"3b",x"5f",x"5f",x"5f",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5f",x"3f",x"3f",x"5f",x"7b",x"97",x"6e",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"8e",x"ff",x"ff",x"f9",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"80",x"84",x"d6",x"df",x"ff",x"ff",x"fa",x"f1",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e8",x"e4",x"e4",x"a4",x"84",x"88",x"d6",x"ff",x"ff",x"fa",x"f5",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"c8",x"a4",x"64",x"b2",x"fb",x"ff",x"ff",x"ff",x"f6",x"e8",x"c4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"a4",x"88",x"b2",x"df",x"ff",x"db",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"49",x"49",x"69",x"69",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"69",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"04",x"24",x"00",x"00",x"00",x"24",x"45",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"92",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"bf",x"7f",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"57",x"52",x"4e",x"2d",x"29",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"6a",x"d7",x"ff",x"fa",x"f5",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"84",x"84",x"ad",x"fb",x"ff",x"df",x"92",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"92",x"fb",x"ff",x"fa",x"f0",x"ec",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"c4",x"80",x"84",x"d6",x"ff",x"ff",x"db",x"db",x"ff",x"ff",x"f6",x"cc",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"c8",x"c8",x"a4",x"80",x"40",x"64",x"8d",x"da",x"ff",x"ff",x"bb",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"09",x"32",x"57",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"5b",x"5b",x"77",x"72",x"6e",x"89",x"84",x"a4",x"89",x"72",x"77",x"77",x"77",x"72",x"89",x"a0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"80",x"60",x"20",x"00",x"00",x"00",x"24",x"24",x"44",x"48",x"49",x"49",x"49",x"29",x"25",x"24",x"04",x"00",x"00",x"00",x"00",x"29",x"96",x"fb",x"fe",x"fa",x"f1",x"d0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"a8",x"84",x"89",x"d7",x"ff",x"ff",x"b6",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"44",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"00",x"00",x"20",x"40",x"60",x"60",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"c0",x"e0",x"c0",x"c0",x"a0",x"a9",x"92",x"76",x"5b",x"7b",x"77",x"92",x"a9",x"a5",x"c4",x"e0",x"e0",x"e0",x"e0",x"c4",x"a5",x"8d",x"92",x"77",x"7b",x"5b",x"5b",x"5b",x"5b",x"5f",x"5f",x"5f",x"5b",x"3b",x"3b",x"5f",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5f",x"5f",x"5b",x"56",x"4e",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"69",x"d7",x"ff",x"fe",x"f9",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e4",x"c4",x"80",x"a9",x"d6",x"ff",x"ff",x"ff",x"f6",x"f1",x"c8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"80",x"84",x"ad",x"db",x"ff",x"ff",x"f5",x"f5",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"a4",x"84",x"89",x"d6",x"ff",x"ff",x"ff",x"fa",x"f1",x"e8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"a4",x"80",x"89",x"d6",x"ff",x"ff",x"b6",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"44",x"49",x"49",x"69",x"69",x"6d",x"6d",x"4d",x"4d",x"4d",x"49",x"49",x"49",x"48",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"29",x"4d",x"72",x"96",x"72",x"29",x"00",x"00",x"24",x"24",x"29",x"49",x"49",x"49",x"6d",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"92",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"9f",x"7b",x"5b",x"5f",x"5f",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5f",x"5b",x"3b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"5b",x"5b",x"7b",x"57",x"57",x"2e",x"29",x"05",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"92",x"fb",x"fb",x"f6",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"c8",x"80",x"84",x"d6",x"ff",x"ff",x"bb",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"b7",x"ff",x"fa",x"f5",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"c4",x"a4",x"84",x"ad",x"fb",x"ff",x"ff",x"b7",x"b7",x"db",x"ff",x"fa",x"d1",x"a8",x"c8",x"c8",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"c8",x"a4",x"a4",x"84",x"84",x"60",x"64",x"b2",x"db",x"ff",x"ff",x"db",x"92",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"09",x"32",x"57",x"7b",x"5b",x"3b",x"37",x"3b",x"5b",x"5b",x"57",x"57",x"72",x"8e",x"85",x"80",x"85",x"89",x"72",x"76",x"57",x"76",x"6e",x"85",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"40",x"20",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"48",x"49",x"45",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"6e",x"db",x"ff",x"fa",x"f5",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"e8",x"e8",x"e8",x"ec",x"c8",x"84",x"84",x"ad",x"fb",x"ff",x"db",x"6d",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"00",x"00",x"20",x"40",x"60",x"60",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a5",x"8e",x"76",x"7b",x"5b",x"77",x"92",x"8d",x"a5",x"c4",x"c4",x"e0",x"e0",x"e0",x"c0",x"c5",x"ad",x"92",x"76",x"7b",x"5b",x"5b",x"5b",x"5b",x"5f",x"5f",x"5f",x"5b",x"3b",x"3b",x"3b",x"3f",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"56",x"2d",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"92",x"fb",x"ff",x"fa",x"f5",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"84",x"88",x"b1",x"da",x"ff",x"ff",x"fb",x"f6",x"ed",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"80",x"89",x"d6",x"ff",x"ff",x"fa",x"f5",x"f0",x"f0",x"f0",x"ec",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"80",x"84",x"ad",x"db",x"ff",x"ff",x"ff",x"f6",x"ed",x"e8",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c8",x"84",x"60",x"b2",x"fb",x"ff",x"db",x"6e",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"44",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"28",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"09",x"2e",x"52",x"56",x"9b",x"bf",x"bb",x"72",x"00",x"00",x"00",x"04",x"24",x"44",x"24",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"6d",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"bf",x"9f",x"7f",x"7f",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5f",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"57",x"32",x"2d",x"05",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6e",x"db",x"ff",x"fa",x"f5",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"ec",x"e8",x"a8",x"84",x"89",x"da",x"ff",x"ff",x"92",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"05",x"72",x"ff",x"ff",x"fa",x"f1",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"c8",x"84",x"8d",x"d6",x"ff",x"ff",x"db",x"4e",x"6e",x"b6",x"ff",x"fb",x"d1",x"a8",x"a8",x"c8",x"e8",x"e8",x"c8",x"e8",x"e8",x"e8",x"e8",x"c8",x"c8",x"a8",x"84",x"64",x"64",x"64",x"64",x"8d",x"d6",x"ff",x"ff",x"ff",x"db",x"92",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"09",x"2e",x"52",x"5b",x"5b",x"37",x"3b",x"3b",x"3b",x"37",x"37",x"77",x"92",x"8e",x"85",x"80",x"85",x"69",x"72",x"56",x"57",x"52",x"6d",x"64",x"80",x"a0",x"a0",x"a0",x"80",x"60",x"60",x"20",x"20",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"44",x"24",x"24",x"24",x"04",x"00",x"00",x"00",x"00",x"49",x"b6",x"ff",x"fa",x"f5",x"f1",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"ec",x"a8",x"64",x"89",x"d6",x"ff",x"ff",x"b6",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"24",x"24",x"00",x"00",x"20",x"40",x"40",x"60",x"60",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"80",x"89",x"72",x"57",x"5b",x"77",x"72",x"8d",x"a4",x"a0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a5",x"a9",x"92",x"7b",x"7b",x"5f",x"5b",x"5b",x"5b",x"5b",x"5f",x"5b",x"5b",x"5b",x"5b",x"3f",x"3f",x"3f",x"5b",x"5b",x"5b",x"5b",x"7f",x"7f",x"7b",x"56",x"09",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"d7",x"ff",x"fa",x"f9",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"a4",x"64",x"ad",x"d6",x"ff",x"ff",x"ff",x"fa",x"ed",x"e8",x"e4",x"e4",x"e8",x"e8",x"e4",x"e4",x"e4",x"c4",x"a4",x"64",x"ad",x"fb",x"ff",x"ff",x"f5",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"60",x"84",x"d6",x"ff",x"ff",x"ff",x"fa",x"f1",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"a4",x"64",x"68",x"d6",x"ff",x"ff",x"92",x"29",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"45",x"45",x"45",x"45",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"05",x"2d",x"52",x"56",x"5b",x"5b",x"7b",x"7b",x"7b",x"bf",x"df",x"bb",x"49",x"00",x"00",x"00",x"04",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"6d",x"6d",x"49",x"24",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"df",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"bf",x"9f",x"bf",x"bf",x"9b",x"97",x"77",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"57",x"57",x"52",x"2e",x"29",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"92",x"fb",x"ff",x"f6",x"f1",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"ec",x"c8",x"84",x"88",x"b1",x"db",x"ff",x"db",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"b7",x"ff",x"fa",x"f5",x"cc",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"a4",x"64",x"b1",x"fb",x"ff",x"db",x"92",x"05",x"29",x"92",x"ff",x"ff",x"fb",x"d1",x"ac",x"88",x"a4",x"84",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"64",x"64",x"89",x"ad",x"b2",x"db",x"ff",x"ff",x"ff",x"ff",x"92",x"49",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"05",x"29",x"52",x"57",x"5b",x"5b",x"3b",x"17",x"17",x"3b",x"5b",x"77",x"92",x"69",x"64",x"60",x"65",x"69",x"52",x"56",x"52",x"4e",x"45",x"60",x"80",x"80",x"80",x"80",x"60",x"40",x"40",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"6e",x"db",x"ff",x"fa",x"f5",x"d0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"c8",x"84",x"64",x"b1",x"fb",x"ff",x"db",x"6e",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"20",x"40",x"40",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"a0",x"80",x"85",x"6e",x"57",x"37",x"57",x"72",x"8d",x"a4",x"a0",x"c0",x"e0",x"e0",x"e0",x"c0",x"a5",x"89",x"92",x"77",x"7b",x"5f",x"5f",x"5b",x"5b",x"7b",x"5f",x"3f",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"5f",x"7f",x"7f",x"7b",x"52",x"29",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"92",x"fb",x"ff",x"fa",x"f5",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e4",x"c4",x"84",x"64",x"b6",x"ff",x"ff",x"ff",x"fb",x"f6",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a4",x"60",x"69",x"b6",x"ff",x"ff",x"fa",x"f5",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"a4",x"60",x"89",x"db",x"ff",x"ff",x"ff",x"f6",x"ed",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c8",x"80",x"64",x"8d",x"ff",x"ff",x"db",x"69",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"29",x"2d",x"4e",x"52",x"77",x"7b",x"7b",x"5f",x"5f",x"7b",x"7b",x"9b",x"bb",x"ff",x"ff",x"b6",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"92",x"92",x"6d",x"49",x"24",x"24",x"6d",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"df",x"ff",x"db",x"d6",x"b2",x"92",x"92",x"92",x"97",x"77",x"77",x"57",x"5b",x"3b",x"3b",x"3b",x"3b",x"57",x"57",x"57",x"32",x"2d",x"05",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"d7",x"ff",x"fa",x"f5",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"a8",x"84",x"ad",x"d6",x"df",x"df",x"b7",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"92",x"db",x"ff",x"fa",x"f1",x"cc",x"ec",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"c4",x"84",x"64",x"b6",x"ff",x"ff",x"b7",x"49",x"00",x"00",x"6e",x"db",x"ff",x"ff",x"fa",x"d2",x"ad",x"89",x"88",x"64",x"64",x"64",x"64",x"64",x"64",x"64",x"68",x"89",x"91",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"49",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"29",x"32",x"57",x"5b",x"37",x"17",x"17",x"37",x"5b",x"57",x"52",x"4e",x"69",x"64",x"60",x"45",x"49",x"2e",x"32",x"32",x"49",x"44",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"04",x"b6",x"ff",x"fb",x"f5",x"f0",x"cc",x"ec",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"a4",x"84",x"88",x"d6",x"ff",x"ff",x"b6",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"20",x"20",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"84",x"69",x"52",x"57",x"37",x"52",x"6d",x"84",x"a4",x"c0",x"c0",x"e0",x"e0",x"c0",x"a5",x"89",x"92",x"77",x"7b",x"5f",x"5f",x"5b",x"5b",x"5b",x"5f",x"3f",x"3b",x"3b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5f",x"5f",x"7b",x"52",x"29",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"29",x"db",x"ff",x"ff",x"f5",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e4",x"a0",x"84",x"89",x"da",x"ff",x"ff",x"ff",x"fa",x"f1",x"c4",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e8",x"a0",x"60",x"92",x"db",x"ff",x"ff",x"fa",x"f1",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"a4",x"84",x"b1",x"ff",x"ff",x"ff",x"fa",x"f1",x"e8",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c8",x"60",x"68",x"b6",x"ff",x"ff",x"b7",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"04",x"04",x"04",x"24",x"24",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"09",x"2d",x"52",x"77",x"7b",x"7b",x"7b",x"7b",x"7b",x"5f",x"5b",x"5b",x"7b",x"9b",x"bb",x"ff",x"ff",x"fb",x"8d",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"6d",x"49",x"24",x"00",x"49",x"b6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"f2",x"cd",x"a9",x"a5",x"a5",x"a9",x"ae",x"8e",x"92",x"77",x"77",x"5b",x"5b",x"57",x"37",x"37",x"37",x"12",x"12",x"32",x"2e",x"29",x"05",x"00",x"00",x"00",x"25",x"6e",x"fb",x"ff",x"f5",x"f1",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"c4",x"84",x"64",x"d6",x"ff",x"ff",x"db",x"6e",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"db",x"ff",x"fa",x"f5",x"f0",x"ec",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"a0",x"84",x"8d",x"db",x"ff",x"ff",x"92",x"25",x"00",x"00",x"01",x"4e",x"b6",x"df",x"ff",x"ff",x"ff",x"fa",x"da",x"d6",x"d6",x"b2",x"b2",x"d2",x"d6",x"d6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"09",x"2e",x"57",x"57",x"37",x"37",x"37",x"33",x"32",x"32",x"32",x"4d",x"48",x"64",x"60",x"45",x"49",x"2e",x"2e",x"2d",x"49",x"44",x"40",x"40",x"60",x"40",x"40",x"40",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"db",x"ff",x"fa",x"f1",x"f0",x"ec",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"c8",x"80",x"64",x"b1",x"ff",x"ff",x"db",x"6e",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"65",x"4e",x"53",x"57",x"52",x"4a",x"65",x"a0",x"c0",x"c0",x"c0",x"e0",x"e0",x"a5",x"89",x"92",x"77",x"5b",x"5f",x"5b",x"5b",x"5b",x"5b",x"5b",x"3f",x"3b",x"3b",x"5b",x"5b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"56",x"2d",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"6e",x"ff",x"ff",x"fa",x"f5",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"80",x"84",x"b2",x"df",x"ff",x"ff",x"fb",x"f2",x"e8",x"e4",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"80",x"64",x"d6",x"ff",x"ff",x"fa",x"f5",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"c4",x"a4",x"84",x"ad",x"da",x"ff",x"ff",x"ff",x"f6",x"ed",x"e4",x"e4",x"e4",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"a4",x"64",x"8d",x"db",x"ff",x"db",x"8e",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"2d",x"2e",x"52",x"57",x"7b",x"7f",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"9b",x"df",x"ff",x"ff",x"ff",x"db",x"8d",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"6d",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"6d",x"6d",x"49",x"00",x"00",x"49",x"92",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"f2",x"e9",x"c4",x"c0",x"c0",x"c0",x"c5",x"c5",x"a5",x"a9",x"8e",x"92",x"72",x"52",x"53",x"57",x"57",x"37",x"32",x"12",x"12",x"0e",x"09",x"09",x"05",x"00",x"00",x"49",x"b6",x"ff",x"fa",x"f5",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"a4",x"84",x"8d",x"da",x"ff",x"ff",x"96",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"6e",x"fb",x"ff",x"f6",x"f0",x"ec",x"ec",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"60",x"84",x"d6",x"ff",x"ff",x"db",x"49",x"00",x"00",x"00",x"00",x"04",x"4d",x"96",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"6e",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"05",x"2e",x"32",x"57",x"57",x"33",x"32",x"32",x"12",x"12",x"31",x"49",x"45",x"60",x"40",x"21",x"25",x"29",x"2d",x"29",x"24",x"20",x"20",x"40",x"40",x"40",x"20",x"20",x"00",x"00",x"00",x"00",x"04",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"92",x"fb",x"ff",x"f6",x"f0",x"ec",x"ec",x"f0",x"f0",x"f0",x"ec",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"c8",x"60",x"88",x"da",x"ff",x"ff",x"b7",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"44",x"49",x"32",x"52",x"52",x"4a",x"65",x"80",x"a0",x"c0",x"c0",x"c0",x"c0",x"a0",x"89",x"92",x"76",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7f",x"7b",x"57",x"32",x"0d",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"96",x"ff",x"ff",x"f5",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"c4",x"80",x"8d",x"da",x"ff",x"ff",x"ff",x"f6",x"ed",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"84",x"89",x"db",x"ff",x"ff",x"f5",x"f1",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"c4",x"c4",x"84",x"64",x"d6",x"ff",x"ff",x"ff",x"fa",x"f1",x"e8",x"e4",x"e4",x"e4",x"e8",x"e8",x"e8",x"e4",x"e8",x"c4",x"80",x"89",x"b6",x"ff",x"ff",x"b7",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"29",x"2d",x"52",x"57",x"57",x"5b",x"5b",x"5f",x"5f",x"5f",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"7b",x"9f",x"df",x"ff",x"ff",x"ff",x"ff",x"b6",x"48",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"6d",x"6d",x"6d",x"24",x"00",x"00",x"49",x"92",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f2",x"ed",x"c9",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a4",x"a9",x"89",x"8d",x"6d",x"6e",x"6e",x"52",x"52",x"32",x"0e",x"0e",x"09",x"09",x"05",x"05",x"00",x"01",x"6e",x"db",x"ff",x"fa",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"c8",x"80",x"84",x"b2",x"fb",x"ff",x"df",x"6e",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"b6",x"ff",x"fb",x"f5",x"cc",x"ec",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"c8",x"a4",x"60",x"8d",x"fb",x"ff",x"df",x"97",x"25",x"00",x"00",x"00",x"00",x"00",x"04",x"49",x"92",x"bb",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"db",x"b7",x"93",x"92",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"05",x"2e",x"52",x"52",x"52",x"32",x"32",x"12",x"12",x"12",x"2d",x"45",x"40",x"40",x"20",x"21",x"05",x"29",x"29",x"04",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"4d",x"db",x"ff",x"fa",x"f5",x"f0",x"ec",x"ec",x"f0",x"f0",x"ec",x"ec",x"ec",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"c8",x"a4",x"64",x"8d",x"ff",x"ff",x"db",x"6e",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"29",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"40",x"20",x"20",x"20",x"44",x"29",x"2e",x"2e",x"4a",x"65",x"60",x"80",x"a0",x"c0",x"a0",x"a0",x"a0",x"85",x"72",x"76",x"57",x"5b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5f",x"7f",x"7f",x"77",x"52",x"09",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"db",x"ff",x"fa",x"f5",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"c4",x"a4",x"84",x"b2",x"ff",x"ff",x"ff",x"fb",x"f1",x"e8",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e8",x"e4",x"c4",x"80",x"84",x"b2",x"ff",x"ff",x"fa",x"f5",x"f0",x"ec",x"ec",x"ec",x"ec",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"c4",x"a4",x"84",x"89",x"fb",x"ff",x"ff",x"ff",x"f6",x"ed",x"e8",x"e4",x"e4",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"a0",x"60",x"ad",x"db",x"ff",x"df",x"92",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"09",x"32",x"56",x"5b",x"7f",x"7f",x"7f",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5f",x"5f",x"5b",x"5b",x"5b",x"7b",x"7f",x"9f",x"bf",x"df",x"ff",x"ff",x"ff",x"ff",x"df",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"49",x"6d",x"92",x"92",x"92",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"6d",x"6d",x"6d",x"49",x"24",x"00",x"00",x"24",x"6d",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"f6",x"f2",x"c9",x"c4",x"c0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"c4",x"c4",x"a4",x"80",x"84",x"65",x"69",x"69",x"49",x"4d",x"2d",x"29",x"09",x"09",x"05",x"00",x"00",x"49",x"b2",x"ff",x"fa",x"f5",x"f0",x"f0",x"ec",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"a4",x"84",x"89",x"fa",x"ff",x"df",x"b7",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"8e",x"fb",x"fb",x"f6",x"f1",x"ec",x"ec",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"a4",x"84",x"88",x"b2",x"ff",x"ff",x"bb",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"6d",x"92",x"96",x"b7",x"db",x"db",x"df",x"df",x"db",x"bb",x"96",x"72",x"49",x"25",x"21",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"05",x"29",x"2e",x"2e",x"2e",x"2e",x"2e",x"0e",x"0a",x"09",x"25",x"20",x"20",x"20",x"00",x"04",x"05",x"05",x"04",x"00",x"00",x"00",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"92",x"ff",x"fa",x"f5",x"f0",x"ec",x"ec",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"a4",x"84",x"89",x"b6",x"ff",x"ff",x"b7",x"29",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"00",x"04",x"25",x"29",x"2e",x"29",x"45",x"60",x"80",x"80",x"a0",x"a0",x"80",x"80",x"85",x"69",x"52",x"57",x"57",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5f",x"7b",x"57",x"4e",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"b6",x"ff",x"fe",x"fa",x"f5",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"a0",x"84",x"ad",x"d6",x"ff",x"ff",x"ff",x"f6",x"ed",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e8",x"e8",x"c4",x"a4",x"60",x"ad",x"db",x"ff",x"fe",x"fa",x"f1",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"a4",x"80",x"88",x"b2",x"ff",x"ff",x"ff",x"fa",x"f2",x"ed",x"e4",x"e4",x"e4",x"e4",x"e4",x"e8",x"e8",x"e8",x"c4",x"80",x"64",x"d6",x"ff",x"ff",x"b7",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"05",x"29",x"2d",x"52",x"56",x"5b",x"5b",x"5b",x"5f",x"7b",x"7b",x"7b",x"7b",x"9b",x"9b",x"9b",x"9b",x"9b",x"bf",x"bf",x"bf",x"9f",x"bf",x"bf",x"bf",x"df",x"df",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"df",x"db",x"ff",x"db",x"db",x"db",x"ff",x"db",x"92",x"49",x"00",x"24",x"49",x"6d",x"92",x"92",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"24",x"24",x"00",x"00",x"24",x"92",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"cd",x"c5",x"c4",x"e0",x"e0",x"e0",x"e0",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"60",x"44",x"44",x"25",x"25",x"25",x"05",x"01",x"00",x"00",x"8e",x"db",x"ff",x"fa",x"f5",x"f0",x"ec",x"ec",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"c4",x"84",x"84",x"ad",x"fb",x"ff",x"db",x"6e",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"b6",x"ff",x"fa",x"f5",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"84",x"60",x"ad",x"db",x"ff",x"ff",x"b2",x"25",x"49",x"29",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"25",x"49",x"49",x"49",x"4e",x"4e",x"4e",x"4a",x"49",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"09",x"09",x"09",x"09",x"05",x"05",x"05",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"4e",x"b7",x"ff",x"fa",x"f5",x"f0",x"ec",x"ec",x"f0",x"f0",x"ec",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"a4",x"64",x"ad",x"db",x"ff",x"ff",x"92",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"29",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"04",x"09",x"09",x"09",x"24",x"40",x"60",x"60",x"80",x"80",x"80",x"80",x"85",x"89",x"72",x"57",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"5b",x"5b",x"7f",x"7b",x"56",x"2d",x"05",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6e",x"db",x"ff",x"fa",x"f5",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"c4",x"80",x"60",x"d2",x"fb",x"ff",x"ff",x"fb",x"f6",x"c8",x"e4",x"e4",x"e4",x"e4",x"e8",x"e4",x"e4",x"e8",x"c4",x"84",x"84",x"b2",x"ff",x"ff",x"fe",x"f5",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"c4",x"a4",x"80",x"89",x"ba",x"ff",x"ff",x"ff",x"f6",x"ed",x"e8",x"e4",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"c8",x"80",x"60",x"89",x"fb",x"ff",x"ff",x"6e",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"09",x"2d",x"52",x"56",x"57",x"5b",x"5b",x"7b",x"7f",x"5f",x"5f",x"7b",x"7b",x"97",x"97",x"92",x"92",x"8e",x"b2",x"d6",x"db",x"ff",x"ff",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"6d",x"24",x"00",x"24",x"6d",x"6d",x"92",x"92",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"92",x"92",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"24",x"92",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f2",x"c9",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"a0",x"80",x"60",x"40",x"40",x"20",x"20",x"20",x"00",x"00",x"00",x"05",x"b7",x"ff",x"ff",x"f5",x"d0",x"f0",x"ec",x"ec",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"c4",x"80",x"89",x"d2",x"ff",x"ff",x"b7",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6e",x"db",x"ff",x"f6",x"f1",x"cc",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"80",x"40",x"d6",x"ff",x"ff",x"db",x"92",x"49",x"92",x"97",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"29",x"92",x"b7",x"6d",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"05",x"05",x"05",x"01",x"25",x"01",x"01",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"21",x"92",x"db",x"ff",x"f6",x"f0",x"ec",x"ec",x"f0",x"f0",x"ec",x"ec",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"c8",x"84",x"64",x"d6",x"ff",x"ff",x"d7",x"6e",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"09",x"09",x"05",x"20",x"40",x"60",x"60",x"60",x"80",x"60",x"60",x"65",x"6e",x"52",x"57",x"57",x"57",x"57",x"57",x"37",x"3b",x"3b",x"3b",x"3b",x"5b",x"5b",x"3b",x"3b",x"3b",x"5b",x"7b",x"7b",x"57",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"b6",x"ff",x"ff",x"f6",x"f5",x"f0",x"f0",x"ec",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"c4",x"80",x"64",x"d6",x"ff",x"ff",x"ff",x"fa",x"f1",x"c8",x"e4",x"e4",x"e4",x"e4",x"e8",x"e8",x"e4",x"e4",x"a0",x"84",x"8d",x"d7",x"ff",x"fe",x"fa",x"f5",x"f0",x"ec",x"ec",x"ec",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"c4",x"a4",x"80",x"ad",x"df",x"ff",x"ff",x"fb",x"f2",x"ed",x"e8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"60",x"64",x"b2",x"ff",x"ff",x"db",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"24",x"2d",x"56",x"57",x"7b",x"7b",x"7f",x"7f",x"5b",x"7b",x"7b",x"7b",x"7b",x"77",x"96",x"92",x"ae",x"aa",x"a5",x"a5",x"a5",x"c9",x"f2",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"b6",x"24",x"00",x"00",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"6d",x"6d",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"04",x"49",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f2",x"ed",x"e4",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"60",x"40",x"40",x"20",x"20",x"00",x"00",x"05",x"4e",x"db",x"ff",x"f6",x"f1",x"f0",x"ec",x"ec",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"e8",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e4",x"a4",x"64",x"b2",x"fb",x"ff",x"db",x"72",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"b6",x"ff",x"ff",x"f5",x"cc",x"cc",x"ec",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"c8",x"84",x"64",x"68",x"db",x"ff",x"ff",x"72",x"4e",x"b6",x"db",x"ff",x"df",x"bb",x"92",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6e",x"db",x"ff",x"ff",x"db",x"b6",x"69",x"21",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"01",x"25",x"29",x"49",x"4e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"69",x"45",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"db",x"ff",x"fa",x"f5",x"f0",x"ec",x"ec",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"80",x"64",x"8d",x"fb",x"ff",x"db",x"6e",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"05",x"00",x"00",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"20",x"25",x"29",x"2a",x"0a",x"2e",x"2e",x"2f",x"4f",x"53",x"53",x"57",x"57",x"5b",x"5b",x"5b",x"1b",x"1b",x"5f",x"7f",x"77",x"52",x"09",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"ff",x"ff",x"fa",x"f5",x"f0",x"ec",x"ec",x"ec",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"80",x"64",x"8d",x"ff",x"ff",x"ff",x"fa",x"f6",x"ed",x"e4",x"e0",x"c0",x"e4",x"e4",x"e4",x"e4",x"e4",x"a4",x"60",x"64",x"d6",x"ff",x"ff",x"fa",x"f5",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"ec",x"ec",x"e8",x"e8",x"e4",x"e4",x"e8",x"a0",x"60",x"ad",x"da",x"ff",x"ff",x"fb",x"f6",x"ed",x"e8",x"e4",x"e4",x"e4",x"e8",x"e8",x"e4",x"e4",x"c4",x"84",x"64",x"91",x"df",x"ff",x"db",x"92",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"29",x"32",x"57",x"5b",x"5b",x"5f",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"97",x"96",x"92",x"92",x"8d",x"a5",x"a5",x"c5",x"c0",x"e0",x"e0",x"c0",x"c0",x"c4",x"cd",x"f2",x"f6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"6d",x"24",x"00",x"00",x"24",x"49",x"4d",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"6d",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"6d",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"d7",x"d2",x"c9",x"c4",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"60",x"60",x"40",x"40",x"20",x"00",x"00",x"29",x"97",x"ff",x"fb",x"f6",x"f1",x"ec",x"ec",x"ec",x"f0",x"ec",x"ec",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"e8",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"c4",x"84",x"68",x"d6",x"ff",x"ff",x"96",x"29",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"db",x"ff",x"fa",x"d1",x"cc",x"cc",x"ec",x"ec",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"60",x"64",x"b1",x"ff",x"ff",x"db",x"4e",x"4e",x"db",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"6e",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"b7",x"ff",x"ff",x"ff",x"ff",x"fb",x"b6",x"8e",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"49",x"6e",x"92",x"b2",x"b6",x"b7",x"ba",x"d6",x"d6",x"db",x"db",x"db",x"d7",x"d7",x"b2",x"92",x"69",x"45",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"6e",x"ff",x"ff",x"f9",x"f0",x"ec",x"ec",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"80",x"84",x"b2",x"ff",x"ff",x"db",x"4a",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"05",x"05",x"09",x"05",x"05",x"05",x"05",x"06",x"0a",x"0a",x"2e",x"2e",x"33",x"57",x"5b",x"5b",x"5b",x"5b",x"56",x"2e",x"05",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"92",x"ff",x"ff",x"f9",x"f0",x"f0",x"ec",x"ec",x"ec",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"60",x"88",x"b6",x"ff",x"ff",x"ff",x"f6",x"ed",x"e8",x"e4",x"e4",x"c4",x"e4",x"e4",x"e4",x"e4",x"c4",x"60",x"64",x"8d",x"fb",x"ff",x"ff",x"f5",x"f1",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"c4",x"80",x"60",x"b2",x"ff",x"ff",x"ff",x"fa",x"f1",x"c8",x"c4",x"e4",x"e4",x"e4",x"e4",x"e8",x"e8",x"e4",x"a0",x"84",x"8d",x"ba",x"df",x"ff",x"b7",x"49",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"29",x"2e",x"52",x"57",x"5b",x"5b",x"5f",x"5f",x"7f",x"7f",x"7b",x"7b",x"97",x"96",x"92",x"b2",x"ad",x"a9",x"a9",x"a5",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c4",x"e9",x"ed",x"f6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"6d",x"24",x"00",x"00",x"00",x"24",x"28",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"d7",x"b2",x"a9",x"a5",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"60",x"60",x"40",x"40",x"20",x"20",x"00",x"00",x"4d",x"db",x"fb",x"fa",x"f5",x"f0",x"ec",x"ec",x"ec",x"f0",x"f0",x"ec",x"ec",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"a4",x"84",x"8d",x"fb",x"ff",x"ff",x"6e",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"92",x"ff",x"ff",x"f6",x"d0",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"a4",x"64",x"89",x"d6",x"ff",x"ff",x"b7",x"72",x"92",x"ff",x"fb",x"f6",x"f1",x"f6",x"fa",x"fb",x"db",x"b2",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6a",x"db",x"ff",x"fa",x"f6",x"f6",x"fa",x"fb",x"fb",x"d7",x"8e",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"49",x"6e",x"b2",x"d6",x"db",x"fb",x"ff",x"ff",x"ff",x"ff",x"fa",x"fa",x"fe",x"ff",x"ff",x"fb",x"ff",x"ff",x"ff",x"fb",x"b2",x"6e",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"b7",x"ff",x"fa",x"f5",x"cc",x"ec",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"a4",x"84",x"ad",x"d6",x"ff",x"df",x"bb",x"6e",x"25",x"25",x"25",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"24",x"25",x"49",x"49",x"49",x"49",x"29",x"25",x"05",x"05",x"01",x"01",x"05",x"0a",x"0e",x"33",x"57",x"7b",x"9b",x"52",x"2d",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6e",x"d7",x"ff",x"fa",x"f5",x"d0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"a4",x"84",x"8d",x"da",x"ff",x"ff",x"fa",x"f1",x"c8",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a4",x"40",x"89",x"d6",x"ff",x"ff",x"fb",x"f5",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"a0",x"60",x"68",x"d6",x"ff",x"ff",x"fb",x"f6",x"ed",x"c4",x"c4",x"e4",x"e8",x"e8",x"e4",x"e8",x"e8",x"c0",x"80",x"64",x"d6",x"ff",x"df",x"df",x"92",x"25",x"00",x"00",x"00",x"00",x"00",x"05",x"2d",x"52",x"57",x"7b",x"7f",x"7f",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"97",x"92",x"b2",x"ae",x"a9",x"c5",x"c5",x"c4",x"c4",x"c4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c9",x"f2",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"ff",x"ff",x"ff",x"df",x"b6",x"24",x"00",x"00",x"00",x"20",x"24",x"24",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"69",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b2",x"8d",x"89",x"a9",x"c5",x"c5",x"e4",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"40",x"40",x"20",x"00",x"00",x"24",x"b2",x"ff",x"fa",x"f5",x"f1",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"80",x"88",x"b6",x"ff",x"ff",x"db",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6e",x"db",x"ff",x"fa",x"f1",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"84",x"84",x"b1",x"ff",x"ff",x"db",x"72",x"72",x"b6",x"ff",x"f6",x"cd",x"cc",x"ed",x"f1",x"fa",x"fa",x"fb",x"da",x"b6",x"6e",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"92",x"ff",x"fb",x"f1",x"cc",x"cc",x"f1",x"f6",x"fa",x"fb",x"fb",x"d7",x"b2",x"6d",x"25",x"00",x"00",x"00",x"00",x"00",x"04",x"6d",x"b2",x"d6",x"fb",x"ff",x"fa",x"fa",x"f6",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"f5",x"d5",x"f5",x"f5",x"f6",x"fa",x"fb",x"fb",x"b2",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"92",x"fb",x"fb",x"f6",x"f1",x"cc",x"ec",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"84",x"a9",x"d2",x"fb",x"ff",x"ff",x"ff",x"db",x"d7",x"d7",x"d7",x"db",x"d7",x"b6",x"92",x"6d",x"45",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"6d",x"92",x"92",x"b6",x"d7",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b7",x"92",x"6e",x"2a",x"05",x"05",x"06",x"4e",x"4e",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"29",x"49",x"4d",x"49",x"21",x"00",x"00",x"00",x"00",x"25",x"92",x"ff",x"fb",x"fa",x"f1",x"d0",x"ec",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"a0",x"80",x"89",x"b6",x"ff",x"ff",x"ff",x"f6",x"e9",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"60",x"44",x"b2",x"ff",x"ff",x"ff",x"fa",x"f1",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"ec",x"ec",x"e8",x"e4",x"e4",x"e4",x"e8",x"c4",x"60",x"64",x"b1",x"ff",x"ff",x"fb",x"f6",x"ed",x"e8",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e8",x"e8",x"80",x"60",x"89",x"fb",x"ff",x"ff",x"b7",x"49",x"00",x"00",x"00",x"29",x"4e",x"73",x"77",x"7b",x"5b",x"5f",x"5f",x"5f",x"5b",x"7b",x"7b",x"7b",x"76",x"92",x"8e",x"89",x"a9",x"a5",x"c5",x"c0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c4",x"a5",x"ad",x"b2",x"bb",x"df",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"6d",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"bb",x"97",x"76",x"92",x"8e",x"ae",x"c9",x"c9",x"c9",x"c5",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"40",x"40",x"20",x"00",x"00",x"00",x"8d",x"db",x"ff",x"f6",x"f1",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"84",x"64",x"8d",x"db",x"ff",x"ff",x"92",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"92",x"ff",x"ff",x"f6",x"f0",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"a4",x"64",x"89",x"d6",x"ff",x"ff",x"b7",x"4e",x"b6",x"fb",x"fb",x"f1",x"cc",x"e8",x"e8",x"ec",x"f1",x"f5",x"fa",x"ff",x"fb",x"d7",x"92",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"db",x"ff",x"fa",x"ed",x"c8",x"c8",x"cc",x"f0",x"f5",x"f6",x"fa",x"fb",x"fb",x"d7",x"92",x"49",x"24",x"04",x"24",x"49",x"6d",x"d6",x"fb",x"fb",x"fa",x"fa",x"f6",x"f5",x"f1",x"d0",x"d0",x"f0",x"f0",x"f0",x"f0",x"f0",x"d0",x"f0",x"f0",x"f0",x"f0",x"f1",x"f5",x"f6",x"fb",x"fb",x"b2",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"b6",x"ff",x"fa",x"f5",x"f1",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"a4",x"84",x"ad",x"f6",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"d6",x"b2",x"6e",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"6d",x"92",x"b6",x"db",x"fb",x"fb",x"fb",x"fb",x"fb",x"fa",x"fa",x"fa",x"fa",x"fa",x"fb",x"ff",x"fb",x"fb",x"b7",x"92",x"4a",x"25",x"05",x"25",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"25",x"45",x"49",x"6d",x"92",x"92",x"b6",x"b7",x"b7",x"25",x"00",x"00",x"00",x"01",x"4e",x"db",x"ff",x"fa",x"f5",x"f0",x"ec",x"ec",x"ec",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"c4",x"80",x"60",x"ad",x"db",x"ff",x"ff",x"f6",x"ed",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"60",x"40",x"8d",x"db",x"ff",x"ff",x"ff",x"f6",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"a4",x"60",x"89",x"d6",x"ff",x"ff",x"f6",x"ed",x"c8",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e8",x"e8",x"a4",x"60",x"89",x"d6",x"ff",x"ff",x"fb",x"6e",x"21",x"00",x"01",x"09",x"32",x"77",x"7b",x"7b",x"7f",x"7f",x"7f",x"7b",x"7b",x"76",x"76",x"92",x"92",x"ad",x"a9",x"a5",x"a4",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"c4",x"c4",x"a5",x"a9",x"a9",x"8d",x"8e",x"92",x"bb",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"92",x"24",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"6d",x"6d",x"49",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"69",x"b6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"9f",x"7f",x"7b",x"7b",x"77",x"96",x"92",x"b2",x"b2",x"ae",x"a9",x"a9",x"a5",x"a5",x"a4",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"60",x"60",x"60",x"40",x"20",x"20",x"00",x"00",x"00",x"b6",x"ff",x"ff",x"f1",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e4",x"e8",x"c4",x"60",x"88",x"b2",x"ff",x"ff",x"bb",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"4d",x"bb",x"ff",x"fa",x"f1",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"80",x"64",x"b1",x"db",x"ff",x"db",x"92",x"6e",x"db",x"ff",x"fa",x"f1",x"e8",x"e8",x"e8",x"e8",x"c8",x"ec",x"f1",x"fa",x"fa",x"fb",x"fb",x"d7",x"92",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"92",x"ff",x"ff",x"f6",x"ec",x"ec",x"e8",x"e8",x"cc",x"ec",x"f1",x"f1",x"f5",x"fa",x"ff",x"fb",x"d7",x"92",x"6e",x"6e",x"b7",x"fb",x"fb",x"f6",x"f2",x"d1",x"cd",x"cc",x"cc",x"ec",x"ec",x"ec",x"ec",x"f0",x"f0",x"f4",x"f0",x"f0",x"f0",x"f4",x"f0",x"f0",x"cc",x"cc",x"f1",x"f6",x"fb",x"fb",x"8e",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"72",x"db",x"ff",x"f6",x"f1",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"a4",x"84",x"cd",x"f6",x"fa",x"fa",x"f6",x"f5",x"f1",x"f1",x"f1",x"f1",x"f5",x"f6",x"f6",x"fa",x"fb",x"fb",x"d7",x"8e",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"49",x"92",x"d6",x"fb",x"fb",x"fb",x"fa",x"fa",x"f6",x"f1",x"f1",x"ed",x"ed",x"ed",x"f1",x"ed",x"cd",x"f1",x"f1",x"f6",x"fa",x"ff",x"ff",x"d7",x"92",x"6a",x"05",x"00",x"00",x"00",x"00",x"05",x"25",x"25",x"49",x"6a",x"92",x"b7",x"d7",x"d6",x"fb",x"fb",x"ff",x"ff",x"ff",x"db",x"49",x"00",x"00",x"00",x"25",x"92",x"ff",x"ff",x"f5",x"f1",x"f0",x"ec",x"ec",x"ec",x"ec",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"c4",x"c4",x"80",x"64",x"d6",x"ff",x"ff",x"f6",x"ed",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"a4",x"40",x"64",x"d6",x"ff",x"ff",x"ff",x"fa",x"f1",x"ec",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"c4",x"a4",x"64",x"b1",x"fb",x"ff",x"fa",x"f1",x"c8",x"c8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"a4",x"60",x"44",x"b2",x"fb",x"ff",x"fb",x"b3",x"25",x"00",x"01",x"0a",x"32",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"9b",x"96",x"92",x"ae",x"ad",x"a9",x"a9",x"c5",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"c5",x"c9",x"a9",x"89",x"8d",x"92",x"92",x"76",x"77",x"9b",x"bf",x"df",x"ff",x"ff",x"ff",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"49",x"04",x"00",x"00",x"20",x"24",x"49",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"92",x"6d",x"6d",x"49",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"92",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"bf",x"7b",x"5b",x"5b",x"5b",x"7b",x"77",x"77",x"7b",x"76",x"76",x"92",x"8e",x"8d",x"89",x"89",x"84",x"a4",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"20",x"20",x"00",x"00",x"29",x"db",x"ff",x"fa",x"f1",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"ec",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"a0",x"60",x"8d",x"da",x"ff",x"ff",x"92",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"92",x"fb",x"ff",x"f1",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e4",x"e8",x"e8",x"a0",x"80",x"88",x"d6",x"ff",x"ff",x"96",x"72",x"92",x"fb",x"ff",x"f5",x"ec",x"e8",x"ec",x"ec",x"ec",x"e8",x"e8",x"ec",x"ec",x"f1",x"f6",x"f6",x"fb",x"fb",x"d7",x"92",x"69",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6e",x"db",x"ff",x"f6",x"f1",x"ec",x"ec",x"e8",x"e8",x"ec",x"ec",x"ec",x"cc",x"cc",x"f1",x"f6",x"fa",x"fb",x"fb",x"db",x"fb",x"fb",x"fb",x"f2",x"ed",x"ed",x"c8",x"c8",x"c8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"f1",x"f1",x"f6",x"ff",x"d7",x"6e",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"b6",x"ff",x"fa",x"f5",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e8",x"e8",x"c8",x"f1",x"f1",x"f1",x"ed",x"cc",x"c8",x"cc",x"cc",x"c8",x"cc",x"cc",x"cc",x"cd",x"f1",x"f2",x"f6",x"fb",x"fb",x"92",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"29",x"6e",x"db",x"fb",x"fb",x"fa",x"f6",x"f5",x"f1",x"ed",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"f0",x"f1",x"f5",x"f6",x"fb",x"fb",x"db",x"92",x"6e",x"6e",x"6e",x"92",x"92",x"b6",x"d7",x"db",x"db",x"fb",x"f7",x"f6",x"d6",x"d6",x"da",x"ff",x"ff",x"ff",x"92",x"25",x"00",x"00",x"00",x"49",x"db",x"ff",x"fa",x"f1",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"c4",x"c4",x"84",x"8d",x"fa",x"fb",x"f6",x"ed",x"c8",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"a0",x"60",x"68",x"92",x"df",x"ff",x"ff",x"fa",x"f5",x"cd",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"a4",x"84",x"8c",x"d6",x"fb",x"f6",x"f2",x"ed",x"c4",x"c4",x"e4",x"e4",x"e4",x"e4",x"e8",x"c4",x"a4",x"60",x"60",x"8d",x"db",x"ff",x"ff",x"b7",x"4a",x"01",x"01",x"05",x"2e",x"57",x"5b",x"7b",x"7b",x"77",x"96",x"92",x"8e",x"a9",x"a9",x"c5",x"c4",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c4",x"c9",x"c9",x"ad",x"8e",x"92",x"92",x"76",x"97",x"9b",x"9b",x"7b",x"7b",x"7b",x"bf",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"92",x"24",x"00",x"00",x"00",x"24",x"24",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"6d",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"24",x"b6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"bf",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"77",x"76",x"96",x"92",x"92",x"8d",x"89",x"84",x"84",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"20",x"00",x"00",x"05",x"6e",x"ff",x"ff",x"f6",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"ec",x"e8",x"e8",x"e8",x"e8",x"e4",x"c4",x"80",x"64",x"b6",x"ff",x"ff",x"bb",x"6d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"db",x"ff",x"fa",x"d1",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e4",x"e8",x"e8",x"80",x"84",x"ad",x"fb",x"ff",x"df",x"72",x"6e",x"db",x"ff",x"fa",x"f1",x"ec",x"e8",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"ed",x"f1",x"f6",x"fa",x"fb",x"fb",x"d6",x"8e",x"69",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"b7",x"ff",x"ff",x"d5",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"cc",x"cc",x"cd",x"f1",x"f6",x"fb",x"fb",x"fb",x"f6",x"f2",x"ed",x"e8",x"e8",x"c8",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"f1",x"fb",x"fb",x"b2",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"db",x"ff",x"fa",x"f1",x"ec",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e8",x"e8",x"ed",x"ed",x"ec",x"e8",x"c8",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c8",x"c8",x"cc",x"f1",x"f6",x"ff",x"db",x"72",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"6d",x"92",x"db",x"ff",x"fb",x"f6",x"f1",x"f1",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"ec",x"cc",x"cc",x"d1",x"f6",x"fa",x"ff",x"fb",x"db",x"b7",x"d6",x"d6",x"fb",x"fb",x"fb",x"fb",x"f6",x"f6",x"f2",x"cd",x"ad",x"b1",x"d6",x"ff",x"ff",x"db",x"49",x"00",x"00",x"00",x"25",x"8e",x"ff",x"ff",x"f6",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"c4",x"c4",x"a8",x"d1",x"f6",x"f6",x"ed",x"e8",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"80",x"64",x"b1",x"db",x"ff",x"ff",x"ff",x"f6",x"d1",x"cc",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"a4",x"84",x"ad",x"f6",x"f6",x"f1",x"ed",x"e8",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e8",x"a4",x"80",x"60",x"89",x"d7",x"ff",x"ff",x"db",x"6e",x"05",x"01",x"05",x"2a",x"52",x"77",x"77",x"96",x"92",x"92",x"ad",x"a9",x"a5",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e0",x"e0",x"c4",x"c4",x"c4",x"c4",x"a9",x"a9",x"a9",x"ae",x"b2",x"96",x"76",x"77",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"7b",x"bf",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f7",x"fb",x"fb",x"ff",x"ff",x"ff",x"db",x"4d",x"00",x"00",x"00",x"24",x"24",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"49",x"49",x"24",x"00",x"00",x"00",x"24",x"6d",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"bf",x"7b",x"5b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"77",x"76",x"72",x"6e",x"69",x"69",x"65",x"60",x"60",x"40",x"40",x"40",x"40",x"20",x"20",x"00",x"00",x"4d",x"bb",x"ff",x"fa",x"f1",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"a0",x"64",x"8d",x"db",x"ff",x"ff",x"92",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"05",x"6e",x"ff",x"ff",x"f6",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e4",x"e8",x"c8",x"60",x"89",x"d6",x"ff",x"ff",x"bb",x"6e",x"92",x"ff",x"ff",x"f6",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"c8",x"c8",x"cc",x"cd",x"f6",x"f6",x"fb",x"fb",x"d6",x"8e",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"db",x"ff",x"fb",x"d1",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"c8",x"c8",x"ed",x"f1",x"f1",x"f1",x"cd",x"c8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"c8",x"cd",x"d6",x"ff",x"db",x"6a",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"92",x"ff",x"ff",x"f5",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e8",x"e8",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"e8",x"e8",x"c8",x"c8",x"cd",x"fb",x"ff",x"db",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"92",x"db",x"ff",x"ff",x"fa",x"f1",x"ed",x"cc",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"ec",x"cc",x"cc",x"f1",x"f5",x"f6",x"fa",x"ff",x"fa",x"fa",x"f6",x"f6",x"f1",x"ed",x"ed",x"e8",x"e8",x"e8",x"84",x"40",x"ad",x"fa",x"ff",x"ff",x"b6",x"24",x"00",x"00",x"00",x"49",x"b6",x"ff",x"fa",x"f1",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"c4",x"cc",x"f1",x"f1",x"ed",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e8",x"c4",x"a0",x"60",x"64",x"8d",x"db",x"ff",x"ff",x"ff",x"fa",x"f1",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e8",x"c4",x"a8",x"f1",x"f1",x"ed",x"c9",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e8",x"a4",x"80",x"64",x"89",x"d2",x"ff",x"ff",x"db",x"72",x"25",x"00",x"05",x"25",x"49",x"92",x"92",x"8e",x"a9",x"c9",x"c9",x"c5",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"c0",x"c0",x"c0",x"a5",x"a9",x"a9",x"ad",x"92",x"96",x"97",x"97",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3f",x"5b",x"5b",x"9f",x"df",x"ff",x"ff",x"ff",x"fb",x"f6",x"ee",x"c9",x"ee",x"f6",x"f6",x"fb",x"ff",x"ff",x"92",x"24",x"00",x"00",x"24",x"29",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"6d",x"6d",x"49",x"49",x"24",x"00",x"00",x"00",x"49",x"b6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"bf",x"7b",x"5b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"5b",x"57",x"77",x"76",x"72",x"6e",x"6d",x"49",x"45",x"44",x"20",x"20",x"20",x"20",x"00",x"00",x"25",x"92",x"ff",x"fb",x"f6",x"f1",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e8",x"c4",x"84",x"88",x"b2",x"ff",x"ff",x"db",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"b7",x"ff",x"fa",x"f1",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"a4",x"64",x"ad",x"fb",x"ff",x"df",x"96",x"92",x"b6",x"ff",x"fa",x"f1",x"cc",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"cd",x"cd",x"d1",x"f6",x"fb",x"fb",x"b7",x"6e",x"25",x"00",x"00",x"00",x"25",x"6e",x"fb",x"fb",x"f6",x"ed",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"ec",x"e8",x"c8",x"c8",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"c8",x"cc",x"b2",x"ff",x"db",x"6e",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6e",x"db",x"ff",x"fa",x"f1",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e8",x"e8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"ec",x"e8",x"e8",x"e8",x"ec",x"e8",x"e8",x"c8",x"c8",x"d2",x"fb",x"ff",x"92",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"69",x"b6",x"fb",x"fb",x"fa",x"f5",x"d1",x"cc",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"f0",x"f1",x"f5",x"f5",x"f1",x"f1",x"f1",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"80",x"40",x"d2",x"ff",x"ff",x"db",x"6e",x"00",x"00",x"00",x"20",x"92",x"fb",x"fb",x"f6",x"f1",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"c4",x"e8",x"ed",x"e8",x"e4",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c8",x"a4",x"60",x"64",x"8d",x"da",x"ff",x"ff",x"ff",x"ff",x"f6",x"f1",x"ec",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e8",x"e8",x"c8",x"ed",x"ed",x"e8",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"c4",x"80",x"60",x"69",x"b2",x"fb",x"ff",x"ff",x"b2",x"25",x"00",x"00",x"00",x"45",x"69",x"a9",x"c9",x"c5",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c5",x"c5",x"a9",x"a9",x"ae",x"92",x"96",x"76",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"3f",x"3b",x"5b",x"bf",x"ff",x"ff",x"ff",x"f6",x"f2",x"e9",x"e5",x"e1",x"c5",x"c9",x"cd",x"f2",x"fb",x"ff",x"db",x"8d",x"00",x"00",x"24",x"49",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"6d",x"6d",x"49",x"49",x"00",x"00",x"00",x"00",x"6d",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"f6",x"f2",x"f6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"bf",x"9b",x"5b",x"5b",x"3f",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"5b",x"57",x"57",x"57",x"52",x"52",x"4e",x"4d",x"29",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"b7",x"ff",x"fa",x"f1",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"a4",x"64",x"8d",x"db",x"ff",x"fb",x"b2",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"92",x"db",x"ff",x"f6",x"f1",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"c4",x"84",x"88",x"d6",x"ff",x"ff",x"bb",x"72",x"b2",x"db",x"ff",x"f6",x"d1",x"c8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"c8",x"a8",x"a8",x"ad",x"d6",x"ff",x"ff",x"db",x"49",x"01",x"00",x"00",x"49",x"b6",x"fb",x"f6",x"f1",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"c4",x"e8",x"c4",x"c4",x"c4",x"e4",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"a8",x"b1",x"ff",x"ff",x"92",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"96",x"ff",x"fb",x"f6",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e8",x"e8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"c8",x"cd",x"f6",x"ff",x"d7",x"6e",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"b6",x"fb",x"ff",x"f6",x"f1",x"ec",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"f0",x"f0",x"ec",x"ec",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"c4",x"c4",x"80",x"64",x"f7",x"ff",x"ff",x"92",x"29",x"00",x"00",x"00",x"49",x"b7",x"ff",x"fa",x"f1",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e8",x"e8",x"e8",x"c8",x"e8",x"e8",x"e4",x"c4",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"84",x"60",x"44",x"8d",x"d6",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"ed",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"a4",x"84",x"60",x"68",x"b2",x"db",x"ff",x"ff",x"b7",x"6d",x"00",x"00",x"20",x"40",x"64",x"a4",x"c4",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c4",x"c4",x"c4",x"a4",x"a5",x"a5",x"a9",x"a9",x"ae",x"92",x"92",x"97",x"7b",x"7b",x"7b",x"5b",x"5f",x"5f",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5f",x"5b",x"7b",x"bf",x"ff",x"ff",x"f6",x"ed",x"e9",x"e4",x"e0",x"e0",x"c0",x"c4",x"c4",x"c9",x"f2",x"f6",x"fb",x"b6",x"20",x"00",x"24",x"49",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"b6",x"92",x"6d",x"49",x"49",x"24",x"00",x"00",x"00",x"24",x"92",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d2",x"ad",x"a9",x"c9",x"ed",x"f2",x"f7",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"9b",x"7b",x"5f",x"5f",x"5b",x"5b",x"5b",x"5b",x"3f",x"3b",x"3b",x"5b",x"5b",x"3b",x"37",x"37",x"17",x"17",x"17",x"12",x"32",x"2e",x"2e",x"2d",x"29",x"05",x"00",x"00",x"00",x"25",x"92",x"db",x"fb",x"f1",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e8",x"c4",x"a4",x"64",x"91",x"ff",x"ff",x"d7",x"8e",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"b7",x"ff",x"fa",x"d1",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"a0",x"60",x"ad",x"db",x"ff",x"df",x"96",x"4d",x"b6",x"fb",x"fb",x"d1",x"cc",x"c8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"a4",x"84",x"84",x"b1",x"ff",x"ff",x"db",x"4e",x"25",x"00",x"21",x"92",x"ff",x"fb",x"f6",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"a4",x"a0",x"a0",x"c4",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"c8",x"a8",x"8d",x"fb",x"ff",x"b7",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"4e",x"db",x"ff",x"f6",x"ed",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"c4",x"c4",x"a4",x"c4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"c8",x"a8",x"d1",x"fb",x"ff",x"92",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"6e",x"d7",x"ff",x"ff",x"f6",x"cd",x"cc",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"c4",x"c4",x"c4",x"c8",x"a4",x"a4",x"c4",x"c4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"ec",x"e8",x"e8",x"e8",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e8",x"e8",x"c4",x"80",x"84",x"ad",x"fb",x"ff",x"df",x"4d",x"00",x"00",x"00",x"25",x"6e",x"db",x"ff",x"f6",x"f1",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e8",x"c8",x"e4",x"e4",x"e4",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"a4",x"40",x"40",x"8d",x"d6",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"f1",x"ec",x"e8",x"e8",x"ec",x"ec",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e8",x"c4",x"80",x"60",x"88",x"b2",x"fb",x"ff",x"ff",x"bb",x"71",x"24",x"00",x"20",x"40",x"60",x"a0",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c4",x"c5",x"a5",x"a9",x"a9",x"ae",x"b2",x"b2",x"b6",x"9b",x"9b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5f",x"5f",x"5b",x"3b",x"5b",x"5b",x"5f",x"7f",x"5b",x"5b",x"7f",x"7b",x"7b",x"bb",x"db",x"f2",x"c9",x"c4",x"e4",x"e0",x"e4",x"e4",x"e4",x"e4",x"c4",x"c4",x"a4",x"a9",x"d2",x"b2",x"20",x"00",x"24",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"ba",x"b6",x"92",x"92",x"6d",x"49",x"49",x"24",x"00",x"00",x"00",x"6d",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"f2",x"ed",x"e9",x"c4",x"c0",x"e0",x"c4",x"c5",x"cd",x"f2",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"bf",x"9b",x"7b",x"5b",x"5f",x"5b",x"3b",x"3b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"3b",x"37",x"37",x"37",x"37",x"33",x"33",x"12",x"0e",x"0e",x"0d",x"09",x"05",x"00",x"00",x"00",x"45",x"db",x"ff",x"fa",x"d1",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e8",x"a4",x"60",x"8d",x"d6",x"ff",x"ff",x"b2",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"92",x"db",x"ff",x"f1",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"80",x"60",x"b6",x"ff",x"ff",x"b7",x"72",x"6e",x"db",x"fb",x"f6",x"f1",x"cc",x"e8",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"a4",x"60",x"88",x"d6",x"ff",x"ff",x"d7",x"29",x"01",x"01",x"49",x"b7",x"ff",x"f6",x"f1",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e8",x"c4",x"a0",x"60",x"64",x"88",x"89",x"ad",x"cd",x"c8",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"c8",x"a4",x"88",x"fa",x"ff",x"db",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"97",x"ff",x"ff",x"f1",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"ec",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"60",x"80",x"60",x"80",x"84",x"c4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"a4",x"cd",x"fa",x"ff",x"b7",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"92",x"db",x"fb",x"fa",x"f5",x"f1",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e8",x"e4",x"c4",x"80",x"60",x"60",x"64",x"84",x"a8",x"c8",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c8",x"a8",x"60",x"89",x"d6",x"ff",x"ff",x"db",x"25",x"00",x"00",x"00",x"29",x"b7",x"ff",x"fa",x"f1",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"80",x"60",x"64",x"8d",x"d6",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"ec",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"e8",x"e8",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"c4",x"80",x"60",x"89",x"b2",x"fb",x"ff",x"ff",x"db",x"4e",x"24",x"00",x"00",x"40",x"60",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c4",x"c4",x"c9",x"a9",x"a9",x"8e",x"92",x"b2",x"97",x"97",x"77",x"7b",x"7b",x"7f",x"5b",x"5b",x"5b",x"5b",x"5f",x"5f",x"5b",x"5b",x"5b",x"5b",x"5b",x"5f",x"5f",x"5b",x"5b",x"7f",x"7b",x"7b",x"7b",x"9b",x"96",x"92",x"b2",x"cd",x"c9",x"c4",x"e0",x"e0",x"e4",x"e4",x"e4",x"c4",x"c4",x"a4",x"80",x"60",x"60",x"64",x"48",x"00",x"00",x"24",x"49",x"6d",x"6d",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"91",x"6d",x"49",x"48",x"24",x"00",x"00",x"00",x"96",x"df",x"ff",x"ff",x"ff",x"fb",x"f6",x"f2",x"ed",x"e5",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c4",x"c9",x"f2",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"bf",x"7f",x"5b",x"5b",x"5b",x"5f",x"5b",x"3b",x"5b",x"5b",x"5b",x"5b",x"3b",x"37",x"3b",x"37",x"37",x"37",x"37",x"33",x"33",x"12",x"0e",x"0e",x"09",x"08",x"05",x"01",x"00",x"21",x"6e",x"ff",x"ff",x"fa",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e8",x"84",x"64",x"b2",x"fb",x"ff",x"db",x"6d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"44",x"d6",x"ff",x"fb",x"cc",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e8",x"e4",x"c4",x"80",x"88",x"da",x"ff",x"ff",x"92",x"6e",x"96",x"ff",x"fb",x"f1",x"ec",x"e8",x"e8",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"ec",x"ec",x"e8",x"ec",x"ec",x"e8",x"e8",x"e4",x"c4",x"84",x"40",x"91",x"db",x"ff",x"fb",x"93",x"01",x"00",x"01",x"8e",x"db",x"ff",x"f2",x"ec",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"c8",x"a4",x"60",x"60",x"69",x"b2",x"b6",x"b6",x"d1",x"cc",x"e8",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"e8",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"c4",x"a4",x"88",x"fa",x"ff",x"db",x"25",x"00",x"01",x"00",x"00",x"00",x"00",x"49",x"db",x"ff",x"fa",x"d0",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"ec",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"80",x"60",x"64",x"69",x"89",x"a9",x"cd",x"ed",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"a4",x"ad",x"d6",x"ff",x"bb",x"6d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"6e",x"db",x"ff",x"fa",x"f1",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e4",x"e8",x"e8",x"e4",x"e8",x"c4",x"a4",x"60",x"40",x"64",x"69",x"8d",x"ad",x"cd",x"cc",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"c4",x"a4",x"64",x"8e",x"db",x"ff",x"df",x"92",x"20",x"00",x"00",x"01",x"6e",x"ff",x"ff",x"f6",x"ec",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"c4",x"84",x"60",x"64",x"ad",x"d6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fa",x"f1",x"e8",x"e8",x"e8",x"ec",x"cc",x"ec",x"ec",x"e8",x"e8",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"c4",x"a4",x"80",x"60",x"65",x"b2",x"fb",x"ff",x"ff",x"db",x"92",x"00",x"00",x"00",x"20",x"60",x"a0",x"c0",x"e0",x"e0",x"e0",x"e5",x"e5",x"c1",x"c0",x"a5",x"a5",x"a9",x"ad",x"ae",x"92",x"92",x"77",x"77",x"9b",x"7b",x"7b",x"5b",x"5b",x"5f",x"5f",x"3b",x"3b",x"5b",x"5b",x"5f",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7f",x"7b",x"7b",x"7b",x"77",x"77",x"96",x"92",x"ae",x"ad",x"a9",x"c5",x"c4",x"c4",x"e0",x"c0",x"c0",x"c4",x"a4",x"a4",x"84",x"80",x"60",x"40",x"20",x"00",x"00",x"00",x"24",x"29",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"96",x"92",x"71",x"6d",x"49",x"49",x"24",x"00",x"00",x"49",x"db",x"ff",x"ff",x"fb",x"f2",x"cd",x"c9",x"c5",x"c4",x"c4",x"e4",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"c4",x"c4",x"c5",x"cd",x"f2",x"fb",x"ff",x"ff",x"df",x"bf",x"9f",x"5b",x"5b",x"5b",x"5f",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"37",x"37",x"33",x"33",x"32",x"0e",x"0e",x"0a",x"09",x"09",x"04",x"00",x"00",x"49",x"b7",x"ff",x"fa",x"f5",x"c8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"a0",x"80",x"89",x"d6",x"ff",x"ff",x"b6",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"6d",x"fb",x"ff",x"fb",x"ec",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e8",x"e8",x"c4",x"60",x"84",x"b2",x"ff",x"ff",x"db",x"6e",x"72",x"db",x"ff",x"fa",x"f1",x"ec",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"a4",x"84",x"68",x"b6",x"ff",x"ff",x"b7",x"4a",x"01",x"00",x"25",x"b7",x"ff",x"fb",x"f1",x"ec",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"a4",x"80",x"84",x"d2",x"fb",x"fb",x"ff",x"fb",x"f6",x"ed",x"e8",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"c8",x"a4",x"88",x"fa",x"ff",x"db",x"25",x"00",x"00",x"00",x"00",x"00",x"25",x"92",x"fb",x"ff",x"f6",x"cc",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"c4",x"a0",x"84",x"ad",x"d6",x"fb",x"fb",x"fb",x"f6",x"ed",x"e8",x"e8",x"e8",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"a4",x"ad",x"d6",x"ff",x"db",x"6e",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"92",x"db",x"fb",x"f6",x"f1",x"cc",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"a4",x"80",x"89",x"b2",x"d6",x"fb",x"fb",x"f6",x"f1",x"ed",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"e8",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"a0",x"60",x"89",x"d2",x"ff",x"ff",x"b6",x"29",x"00",x"00",x"00",x"49",x"b7",x"ff",x"fb",x"f1",x"ec",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"a4",x"80",x"60",x"64",x"ad",x"d6",x"ff",x"ff",x"ff",x"db",x"db",x"ff",x"fb",x"f6",x"ed",x"ec",x"ec",x"e8",x"e8",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e8",x"c8",x"80",x"60",x"60",x"8d",x"b2",x"db",x"ff",x"ff",x"db",x"6d",x"20",x"00",x"00",x"40",x"80",x"a0",x"e0",x"e0",x"e0",x"e0",x"c4",x"c5",x"c5",x"a9",x"89",x"8d",x"92",x"b2",x"96",x"9b",x"9b",x"7b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"3b",x"5b",x"5b",x"5f",x"5b",x"5b",x"5b",x"7f",x"5b",x"5b",x"5b",x"7b",x"9b",x"97",x"b2",x"b2",x"ae",x"a9",x"a9",x"c9",x"c5",x"c5",x"c5",x"c5",x"c4",x"a4",x"a4",x"80",x"60",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"24",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"49",x"24",x"20",x"00",x"24",x"8d",x"ff",x"ff",x"f6",x"d2",x"cd",x"c5",x"c0",x"c0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"c0",x"c4",x"c9",x"d2",x"f6",x"ff",x"ff",x"df",x"9f",x"7b",x"5b",x"5b",x"5f",x"5f",x"5b",x"5b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"3b",x"37",x"37",x"13",x"12",x"12",x"0e",x"0e",x"09",x"09",x"05",x"00",x"00",x"01",x"8e",x"fb",x"fb",x"f6",x"f1",x"c8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e8",x"c4",x"80",x"84",x"ad",x"fb",x"ff",x"df",x"6d",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"b2",x"fb",x"fb",x"f6",x"ec",x"e8",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e8",x"e4",x"a4",x"40",x"8d",x"da",x"ff",x"ff",x"b7",x"6e",x"96",x"ff",x"fb",x"f6",x"ec",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"80",x"84",x"8d",x"da",x"ff",x"ff",x"8e",x"25",x"00",x"01",x"6e",x"ff",x"ff",x"f6",x"f1",x"ec",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"c4",x"80",x"84",x"ad",x"fb",x"ff",x"ff",x"ff",x"ff",x"fa",x"ed",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"a4",x"89",x"fa",x"ff",x"db",x"49",x"00",x"00",x"00",x"00",x"00",x"49",x"b7",x"ff",x"fa",x"f5",x"cc",x"c8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"c4",x"a4",x"80",x"a9",x"d6",x"fb",x"ff",x"ff",x"ff",x"fa",x"f1",x"ec",x"e8",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"a4",x"a9",x"d6",x"ff",x"db",x"6e",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"92",x"db",x"ff",x"f6",x"f1",x"cd",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e8",x"c4",x"84",x"64",x"b1",x"fb",x"ff",x"ff",x"ff",x"fa",x"f6",x"ed",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e4",x"c4",x"80",x"40",x"b2",x"fb",x"ff",x"df",x"72",x"00",x"00",x"00",x"00",x"6e",x"db",x"ff",x"fa",x"f1",x"ec",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"80",x"60",x"60",x"88",x"b1",x"d6",x"ff",x"ff",x"db",x"b7",x"b7",x"db",x"ff",x"fb",x"d1",x"cc",x"e8",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"80",x"60",x"64",x"8d",x"d6",x"ff",x"ff",x"ff",x"db",x"8e",x"44",x"00",x"00",x"20",x"40",x"80",x"a0",x"c0",x"c0",x"c5",x"a9",x"a9",x"ad",x"ad",x"92",x"96",x"96",x"97",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5f",x"5f",x"5f",x"3f",x"3b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"77",x"76",x"72",x"92",x"92",x"ae",x"ad",x"c9",x"c9",x"c5",x"c5",x"c5",x"a1",x"a0",x"a0",x"80",x"80",x"60",x"60",x"40",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"69",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"92",x"92",x"6d",x"4d",x"24",x"00",x"00",x"69",x"d6",x"fb",x"d2",x"cd",x"c9",x"c5",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e4",x"e0",x"e0",x"c0",x"c0",x"c9",x"cd",x"f6",x"fb",x"df",x"bb",x"9b",x"7b",x"5b",x"5f",x"5f",x"5b",x"5b",x"3b",x"3b",x"37",x"3b",x"3b",x"3b",x"3b",x"37",x"17",x"13",x"12",x"0e",x"0e",x"09",x"09",x"05",x"00",x"00",x"00",x"29",x"b7",x"ff",x"fb",x"f1",x"ec",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"c4",x"80",x"89",x"d6",x"ff",x"ff",x"b7",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6e",x"d7",x"fb",x"f6",x"f1",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e8",x"a4",x"60",x"68",x"b6",x"ff",x"ff",x"bb",x"6e",x"72",x"bb",x"ff",x"fa",x"f1",x"c8",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"80",x"84",x"b2",x"ff",x"ff",x"db",x"4a",x"00",x"00",x"29",x"92",x"ff",x"fb",x"f1",x"ed",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"a4",x"60",x"89",x"d6",x"ff",x"ff",x"ff",x"ff",x"ff",x"f6",x"ec",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e8",x"c4",x"84",x"89",x"fb",x"ff",x"db",x"45",x"00",x"00",x"00",x"00",x"00",x"92",x"ff",x"fb",x"f6",x"f1",x"cc",x"e8",x"e8",x"ec",x"ec",x"ec",x"e8",x"e8",x"ec",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"80",x"84",x"b1",x"fb",x"ff",x"ff",x"ff",x"ff",x"fa",x"f1",x"ec",x"e8",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"80",x"a9",x"d6",x"ff",x"db",x"6d",x"20",x"00",x"00",x"00",x"00",x"00",x"25",x"6e",x"db",x"ff",x"fa",x"f1",x"cd",x"cc",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"c8",x"84",x"64",x"89",x"d6",x"ff",x"ff",x"ff",x"ff",x"ff",x"f6",x"ed",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"e8",x"ec",x"e8",x"e4",x"e4",x"e4",x"e4",x"a4",x"60",x"64",x"fa",x"ff",x"ff",x"b7",x"49",x"00",x"00",x"00",x"05",x"b6",x"ff",x"fb",x"f6",x"f1",x"e8",x"e8",x"e8",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"80",x"40",x"44",x"89",x"b6",x"db",x"ff",x"ff",x"db",x"92",x"6e",x"92",x"fb",x"ff",x"f6",x"cd",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"c4",x"c4",x"80",x"40",x"64",x"8d",x"da",x"ff",x"ff",x"ff",x"bb",x"8e",x"24",x"20",x"00",x"20",x"40",x"60",x"80",x"a0",x"a5",x"a9",x"8d",x"92",x"92",x"96",x"96",x"9b",x"7b",x"7b",x"7b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5f",x"5f",x"5f",x"5f",x"5f",x"5b",x"7b",x"7b",x"97",x"97",x"97",x"b7",x"b7",x"92",x"92",x"8d",x"89",x"a9",x"a5",x"a5",x"a5",x"a5",x"a4",x"84",x"84",x"80",x"80",x"60",x"60",x"40",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"24",x"24",x"24",x"49",x"49",x"6d",x"8e",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"92",x"92",x"6d",x"49",x"24",x"00",x"00",x"69",x"b2",x"8d",x"89",x"a4",x"c4",x"c4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c4",x"c4",x"c4",x"c9",x"d2",x"b7",x"97",x"97",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"37",x"37",x"37",x"37",x"17",x"13",x"12",x"12",x"0e",x"0a",x"09",x"05",x"05",x"00",x"00",x"05",x"72",x"db",x"ff",x"f6",x"ed",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"c4",x"a4",x"84",x"b2",x"fb",x"ff",x"db",x"6e",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"b7",x"ff",x"fb",x"f1",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e8",x"e8",x"e8",x"c4",x"80",x"60",x"91",x"db",x"ff",x"ff",x"92",x"49",x"b7",x"ff",x"fb",x"f1",x"cc",x"e8",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"c4",x"84",x"8d",x"d6",x"ff",x"df",x"92",x"25",x"00",x"01",x"6e",x"db",x"ff",x"f6",x"ed",x"ec",x"e8",x"e8",x"ec",x"ec",x"ec",x"e8",x"e8",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"c4",x"84",x"84",x"b1",x"fb",x"ff",x"ff",x"ff",x"ff",x"fa",x"f1",x"c8",x"c8",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e8",x"a0",x"84",x"ad",x"fb",x"ff",x"b7",x"25",x"00",x"00",x"00",x"00",x"29",x"bb",x"ff",x"fa",x"f1",x"cc",x"c8",x"e8",x"e8",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"80",x"60",x"ad",x"d6",x"ff",x"ff",x"ff",x"ff",x"ff",x"f6",x"cc",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"80",x"a9",x"f6",x"ff",x"db",x"6d",x"20",x"00",x"00",x"00",x"00",x"04",x"6e",x"db",x"ff",x"fa",x"f1",x"ec",x"ec",x"e8",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"c4",x"60",x"64",x"d2",x"ff",x"ff",x"df",x"df",x"ff",x"fa",x"f1",x"cc",x"e8",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"ec",x"e8",x"e4",x"e4",x"e4",x"c4",x"80",x"64",x"8d",x"ff",x"ff",x"ff",x"6e",x"24",x"00",x"00",x"00",x"4d",x"db",x"ff",x"f6",x"f1",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"c4",x"a0",x"80",x"60",x"40",x"89",x"b2",x"db",x"ff",x"ff",x"ff",x"bb",x"6e",x"05",x"4a",x"b6",x"ff",x"fa",x"f5",x"cc",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e8",x"e4",x"e4",x"e4",x"c4",x"c4",x"a4",x"60",x"40",x"64",x"8d",x"d6",x"ff",x"ff",x"ff",x"df",x"92",x"29",x"00",x"00",x"00",x"00",x"20",x"44",x"69",x"8e",x"b2",x"b2",x"96",x"77",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"3b",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"9b",x"97",x"93",x"8e",x"8e",x"89",x"89",x"89",x"a8",x"a8",x"a4",x"a4",x"a4",x"a4",x"a4",x"80",x"60",x"40",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"24",x"28",x"29",x"29",x"49",x"49",x"6d",x"8d",x"92",x"b2",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"d7",x"b6",x"92",x"92",x"6d",x"49",x"24",x"00",x"00",x"44",x"69",x"44",x"60",x"80",x"a0",x"a0",x"c4",x"c4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c9",x"ce",x"ae",x"92",x"92",x"96",x"77",x"77",x"7b",x"7b",x"7b",x"57",x"57",x"37",x"37",x"37",x"37",x"13",x"12",x"0e",x"0e",x"09",x"05",x"05",x"00",x"00",x"00",x"25",x"97",x"ff",x"ff",x"f1",x"ec",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"a0",x"80",x"89",x"d6",x"ff",x"ff",x"b7",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6e",x"db",x"ff",x"f6",x"ed",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e8",x"e4",x"a0",x"60",x"68",x"db",x"ff",x"ff",x"bb",x"6e",x"4d",x"db",x"ff",x"f6",x"cd",x"c8",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"a0",x"89",x"b2",x"ff",x"ff",x"db",x"49",x"01",x"00",x"25",x"b6",x"ff",x"fb",x"f1",x"ec",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"ec",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"80",x"89",x"d6",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"ed",x"c8",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e8",x"80",x"84",x"b2",x"ff",x"ff",x"b6",x"24",x"00",x"00",x"00",x"04",x"72",x"df",x"ff",x"f5",x"ec",x"c8",x"e8",x"e8",x"e8",x"e8",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"80",x"64",x"d2",x"ff",x"ff",x"df",x"ff",x"ff",x"fa",x"f1",x"c8",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e8",x"c8",x"80",x"ad",x"fa",x"ff",x"db",x"69",x"00",x"00",x"00",x"00",x"00",x"4d",x"b6",x"ff",x"fb",x"f5",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e8",x"e4",x"a4",x"60",x"89",x"fb",x"ff",x"ff",x"df",x"ff",x"ff",x"f6",x"cd",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"c4",x"80",x"88",x"b2",x"ff",x"ff",x"db",x"25",x"00",x"00",x"00",x"25",x"96",x"ff",x"fb",x"f1",x"cc",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"a0",x"60",x"60",x"64",x"89",x"d6",x"fb",x"ff",x"ff",x"ff",x"bb",x"6e",x"05",x"01",x"6e",x"db",x"fb",x"f6",x"d1",x"cc",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"a0",x"80",x"60",x"64",x"69",x"92",x"db",x"ff",x"ff",x"ff",x"db",x"92",x"29",x"00",x"00",x"00",x"00",x"25",x"49",x"6d",x"72",x"97",x"9b",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5f",x"5f",x"5f",x"3b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"7b",x"97",x"77",x"77",x"96",x"92",x"b2",x"ad",x"a9",x"a5",x"a4",x"84",x"84",x"a0",x"a0",x"80",x"80",x"60",x"60",x"40",x"40",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"24",x"24",x"24",x"29",x"29",x"49",x"49",x"49",x"4d",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"d7",x"b6",x"92",x"92",x"6d",x"4d",x"49",x"24",x"00",x"00",x"20",x"20",x"40",x"60",x"60",x"60",x"80",x"84",x"84",x"a4",x"a4",x"c4",x"c4",x"e4",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"c5",x"c5",x"a9",x"a9",x"8d",x"8e",x"92",x"92",x"92",x"96",x"72",x"77",x"57",x"57",x"57",x"33",x"32",x"32",x"0e",x"0e",x"09",x"05",x"05",x"00",x"00",x"00",x"4d",x"df",x"ff",x"fa",x"f1",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"80",x"60",x"b1",x"db",x"ff",x"df",x"92",x"05",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"b7",x"ff",x"ff",x"f1",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"c4",x"60",x"64",x"91",x"ff",x"ff",x"db",x"72",x"4e",x"72",x"ff",x"ff",x"f1",x"c8",x"c8",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c8",x"a0",x"80",x"ad",x"db",x"ff",x"ff",x"97",x"25",x"00",x"01",x"6e",x"db",x"ff",x"f6",x"ed",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"c4",x"80",x"60",x"b2",x"fb",x"ff",x"ff",x"ff",x"ff",x"fa",x"f1",x"ec",x"c8",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"c4",x"60",x"88",x"d6",x"ff",x"ff",x"92",x"24",x"00",x"00",x"00",x"25",x"b7",x"ff",x"fb",x"f1",x"e8",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"84",x"89",x"fb",x"ff",x"ff",x"db",x"ff",x"ff",x"f6",x"d1",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"a4",x"84",x"ad",x"fb",x"ff",x"d7",x"49",x"00",x"00",x"00",x"00",x"25",x"b6",x"fb",x"fb",x"f6",x"ed",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e8",x"c4",x"80",x"84",x"b2",x"ff",x"ff",x"df",x"ff",x"ff",x"ff",x"d1",x"cc",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"a4",x"64",x"ad",x"db",x"ff",x"df",x"92",x"00",x"00",x"00",x"00",x"4d",x"db",x"ff",x"fa",x"ed",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e0",x"e4",x"e4",x"c8",x"c4",x"80",x"60",x"44",x"64",x"ae",x"d7",x"ff",x"ff",x"ff",x"ff",x"b7",x"6e",x"00",x"00",x"25",x"b7",x"ff",x"fa",x"f1",x"cc",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"c4",x"c4",x"c4",x"a0",x"60",x"40",x"64",x"8d",x"b6",x"ff",x"ff",x"ff",x"ff",x"fb",x"92",x"49",x"00",x"00",x"00",x"00",x"29",x"4e",x"92",x"97",x"7b",x"7b",x"5b",x"5b",x"3b",x"5b",x"5b",x"5b",x"5f",x"5b",x"3f",x"3f",x"3f",x"5f",x"5b",x"5b",x"5b",x"7b",x"7b",x"9b",x"97",x"96",x"b6",x"b2",x"ae",x"ad",x"a9",x"a9",x"a9",x"a4",x"a4",x"c4",x"c8",x"a8",x"a4",x"80",x"60",x"60",x"40",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"24",x"24",x"24",x"24",x"24",x"28",x"28",x"29",x"49",x"49",x"49",x"4d",x"4d",x"6d",x"6d",x"72",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"72",x"6d",x"49",x"24",x"20",x"00",x"00",x"20",x"20",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"40",x"60",x"80",x"80",x"a0",x"a4",x"a4",x"c4",x"c4",x"e4",x"e4",x"e0",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c5",x"a5",x"a5",x"a5",x"85",x"89",x"89",x"8d",x"6e",x"6e",x"4e",x"4e",x"4e",x"2e",x"2e",x"2e",x"09",x"09",x"05",x"05",x"00",x"00",x"25",x"92",x"ff",x"ff",x"f6",x"cc",x"e8",x"e8",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"80",x"64",x"d6",x"ff",x"ff",x"b7",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"8e",x"fb",x"fb",x"f6",x"cd",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e8",x"e8",x"e4",x"a0",x"80",x"60",x"8d",x"d7",x"ff",x"ff",x"b7",x"49",x"6e",x"bb",x"ff",x"fa",x"f1",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e8",x"e8",x"c4",x"80",x"60",x"b2",x"ff",x"ff",x"bb",x"6e",x"01",x"00",x"25",x"b6",x"fb",x"fb",x"f1",x"ec",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"a4",x"60",x"64",x"d6",x"ff",x"ff",x"df",x"ff",x"fb",x"f6",x"ed",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"c4",x"60",x"89",x"d6",x"ff",x"db",x"92",x"24",x"00",x"00",x"00",x"6e",x"fb",x"ff",x"f6",x"ec",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"60",x"84",x"b2",x"ff",x"ff",x"ff",x"db",x"fb",x"fa",x"f1",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"c4",x"a4",x"88",x"b2",x"ff",x"ff",x"b6",x"45",x"00",x"00",x"00",x"25",x"92",x"ff",x"fb",x"f6",x"d1",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"a4",x"80",x"ad",x"d6",x"ff",x"ff",x"db",x"fb",x"fb",x"f6",x"cd",x"c8",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e8",x"e8",x"a4",x"80",x"88",x"b2",x"ff",x"ff",x"bb",x"49",x"00",x"00",x"00",x"29",x"92",x"ff",x"fa",x"f1",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e8",x"e4",x"c4",x"80",x"60",x"60",x"64",x"89",x"b2",x"d7",x"fb",x"ff",x"ff",x"ff",x"db",x"6e",x"25",x"20",x"00",x"21",x"6e",x"db",x"ff",x"f6",x"ed",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"a4",x"80",x"60",x"60",x"68",x"ad",x"d6",x"fb",x"ff",x"ff",x"ff",x"ff",x"b7",x"6e",x"25",x"00",x"00",x"00",x"05",x"2e",x"56",x"7b",x"7b",x"5b",x"5b",x"3f",x"3f",x"3f",x"5b",x"5f",x"5f",x"5f",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"97",x"96",x"b2",x"ae",x"ad",x"a9",x"a9",x"c9",x"a4",x"c4",x"c4",x"c4",x"c0",x"c0",x"c4",x"e9",x"f2",x"f6",x"ad",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"20",x"24",x"24",x"24",x"44",x"44",x"45",x"49",x"49",x"49",x"49",x"49",x"69",x"6d",x"6d",x"6d",x"6d",x"6e",x"92",x"92",x"b6",x"b6",x"ba",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"40",x"40",x"60",x"64",x"84",x"84",x"a4",x"a0",x"c0",x"c4",x"c4",x"c4",x"c4",x"c4",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a4",x"a4",x"a5",x"85",x"69",x"69",x"69",x"49",x"29",x"29",x"29",x"09",x"05",x"05",x"00",x"00",x"00",x"6e",x"bb",x"ff",x"fa",x"f1",x"c8",x"e8",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"80",x"64",x"8d",x"fb",x"ff",x"df",x"6e",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"44",x"92",x"d7",x"fb",x"f6",x"f1",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e8",x"e8",x"c4",x"80",x"60",x"89",x"b6",x"ff",x"ff",x"db",x"8e",x"25",x"92",x"ff",x"fa",x"f6",x"ed",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"a4",x"60",x"88",x"db",x"ff",x"ff",x"92",x"25",x"01",x"01",x"4a",x"db",x"ff",x"f6",x"cd",x"c8",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"c4",x"a0",x"60",x"89",x"fb",x"ff",x"df",x"ff",x"ff",x"fa",x"f1",x"e8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"c4",x"a4",x"64",x"8d",x"db",x"ff",x"db",x"49",x"00",x"00",x"00",x"49",x"92",x"fb",x"fb",x"f1",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"c4",x"a4",x"60",x"8d",x"d6",x"ff",x"ff",x"ff",x"fb",x"fb",x"f6",x"cd",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"a0",x"80",x"ad",x"d6",x"ff",x"ff",x"92",x"20",x"00",x"00",x"00",x"6d",x"d6",x"ff",x"fa",x"f1",x"cc",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"80",x"64",x"b2",x"ff",x"ff",x"ff",x"ff",x"fb",x"fa",x"f1",x"c8",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"80",x"60",x"ad",x"d7",x"ff",x"ff",x"92",x"05",x"00",x"00",x"00",x"6e",x"db",x"ff",x"f6",x"f1",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"a4",x"80",x"64",x"64",x"6d",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"df",x"b7",x"6e",x"25",x"00",x"00",x"00",x"45",x"97",x"fb",x"fb",x"f1",x"ec",x"e8",x"e8",x"e8",x"e8",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"a0",x"a0",x"80",x"84",x"64",x"68",x"8d",x"b2",x"db",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"49",x"21",x"00",x"00",x"01",x"05",x"2e",x"57",x"5b",x"5b",x"5b",x"3b",x"3f",x"3f",x"3f",x"5f",x"5b",x"7b",x"7b",x"7b",x"7b",x"7b",x"7b",x"97",x"97",x"96",x"92",x"92",x"ae",x"ad",x"a9",x"a9",x"a5",x"a4",x"a0",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e4",x"ed",x"f2",x"fb",x"d6",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"25",x"45",x"45",x"49",x"69",x"69",x"69",x"69",x"69",x"6d",x"6d",x"6d",x"8e",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"ba",x"b6",x"92",x"92",x"92",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"40",x"40",x"60",x"60",x"80",x"80",x"84",x"a4",x"a4",x"c4",x"c4",x"c4",x"c0",x"c0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"60",x"60",x"40",x"20",x"20",x"20",x"04",x"00",x"00",x"00",x"00",x"25",x"b6",x"ff",x"fb",x"f5",x"cc",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"60",x"88",x"d6",x"ff",x"ff",x"bb",x"29",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"8e",x"fb",x"ff",x"fa",x"f1",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"a4",x"60",x"64",x"b6",x"ff",x"ff",x"fb",x"92",x"49",x"4a",x"b7",x"ff",x"f6",x"ed",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"c4",x"80",x"64",x"b1",x"ff",x"ff",x"db",x"49",x"00",x"00",x"25",x"92",x"ff",x"fb",x"f5",x"c8",x"c8",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"c4",x"80",x"85",x"b2",x"ff",x"ff",x"df",x"ff",x"ff",x"f6",x"ed",x"e8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"c0",x"80",x"89",x"d6",x"ff",x"ff",x"b7",x"25",x"00",x"00",x"00",x"6e",x"db",x"fb",x"f6",x"ed",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"c4",x"80",x"64",x"b2",x"fb",x"ff",x"ff",x"ff",x"ff",x"fa",x"f1",x"e8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"a0",x"60",x"b1",x"fb",x"ff",x"db",x"4e",x"00",x"00",x"01",x"25",x"b7",x"ff",x"fa",x"f1",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"60",x"88",x"d6",x"ff",x"df",x"ff",x"ff",x"fb",x"f6",x"ed",x"c4",x"c4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"80",x"64",x"d2",x"fb",x"ff",x"db",x"6e",x"00",x"00",x"00",x"21",x"b2",x"ff",x"ff",x"f6",x"ed",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a4",x"80",x"40",x"44",x"8d",x"b6",x"db",x"df",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"49",x"00",x"00",x"00",x"00",x"00",x"69",x"db",x"fb",x"f6",x"ed",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"a0",x"60",x"60",x"60",x"89",x"8d",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"fb",x"b7",x"4d",x"00",x"00",x"00",x"01",x"05",x"0a",x"32",x"57",x"7b",x"5b",x"5b",x"3b",x"3f",x"5f",x"5f",x"7f",x"7b",x"7b",x"77",x"77",x"97",x"97",x"97",x"b6",x"b2",x"ae",x"ad",x"a9",x"a9",x"a5",x"a5",x"a4",x"a4",x"a4",x"a4",x"a0",x"a0",x"a0",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e9",x"f2",x"fb",x"db",x"72",x"29",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"24",x"24",x"24",x"25",x"49",x"49",x"69",x"69",x"69",x"6d",x"6d",x"6d",x"8d",x"8d",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"b6",x"92",x"92",x"92",x"8d",x"6d",x"49",x"49",x"29",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"40",x"40",x"60",x"80",x"80",x"a4",x"a0",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"60",x"40",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"4d",x"db",x"ff",x"f6",x"ed",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"c4",x"a4",x"60",x"ad",x"fb",x"ff",x"db",x"92",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"92",x"db",x"fb",x"f6",x"f1",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"40",x"68",x"b6",x"ff",x"ff",x"ff",x"b7",x"49",x"01",x"93",x"db",x"ff",x"d6",x"cc",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"60",x"89",x"da",x"ff",x"ff",x"b7",x"25",x"00",x"00",x"6a",x"d7",x"ff",x"fa",x"f1",x"c8",x"c8",x"e8",x"e8",x"e8",x"e8",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"a4",x"60",x"a9",x"f7",x"ff",x"ff",x"df",x"ff",x"fa",x"f1",x"e8",x"e4",x"e4",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e8",x"e8",x"e4",x"e8",x"e8",x"e4",x"e4",x"a0",x"60",x"ad",x"db",x"ff",x"df",x"92",x"05",x"00",x"00",x"25",x"b7",x"ff",x"fb",x"f1",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"a0",x"60",x"89",x"d6",x"ff",x"ff",x"ff",x"ff",x"ff",x"f6",x"ed",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"80",x"60",x"d6",x"ff",x"ff",x"b7",x"49",x"00",x"00",x"25",x"92",x"fb",x"ff",x"f6",x"cc",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"c4",x"80",x"64",x"ad",x"db",x"ff",x"df",x"df",x"ff",x"fa",x"f2",x"ed",x"c4",x"e4",x"e8",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e8",x"e4",x"c4",x"a0",x"80",x"89",x"fb",x"ff",x"ff",x"92",x"29",x"00",x"00",x"20",x"69",x"db",x"ff",x"fb",x"d1",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"a0",x"84",x"88",x"ad",x"d6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"45",x"92",x"ff",x"ff",x"f6",x"cc",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"a4",x"80",x"64",x"89",x"b2",x"d6",x"fb",x"ff",x"ff",x"ff",x"ff",x"db",x"b2",x"49",x"25",x"00",x"00",x"00",x"00",x"05",x"2e",x"57",x"57",x"5b",x"5b",x"5b",x"5f",x"5b",x"5f",x"7f",x"9b",x"9b",x"9b",x"96",x"92",x"92",x"8e",x"ad",x"a9",x"a9",x"a9",x"a5",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"85",x"89",x"89",x"89",x"89",x"a5",x"a4",x"c0",x"e0",x"e4",x"e4",x"c0",x"c4",x"c9",x"f6",x"ff",x"db",x"4d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"24",x"25",x"48",x"48",x"49",x"4d",x"4d",x"6d",x"6d",x"71",x"72",x"92",x"92",x"92",x"92",x"92",x"96",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b2",x"92",x"92",x"6d",x"6d",x"4d",x"4d",x"49",x"49",x"49",x"45",x"45",x"44",x"44",x"24",x"24",x"24",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"40",x"40",x"60",x"60",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"60",x"40",x"40",x"20",x"20",x"00",x"00",x"00",x"24",x"92",x"ff",x"ff",x"f2",x"c8",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"84",x"84",x"d2",x"ff",x"ff",x"b7",x"49",x"00",x"00",x"00",x"00",x"25",x"69",x"b2",x"fb",x"fb",x"f6",x"f1",x"c8",x"e4",x"e4",x"e4",x"e8",x"e8",x"e4",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"60",x"64",x"b2",x"ff",x"ff",x"ff",x"db",x"6e",x"01",x"01",x"db",x"ff",x"fa",x"d1",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"c4",x"a0",x"60",x"ad",x"ff",x"ff",x"db",x"6e",x"05",x"00",x"05",x"92",x"fb",x"fb",x"f6",x"ed",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"a0",x"64",x"b2",x"ff",x"ff",x"ff",x"ff",x"ff",x"f6",x"ed",x"e8",x"e4",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e8",x"e4",x"e4",x"e8",x"e8",x"e4",x"c4",x"80",x"60",x"b2",x"ff",x"ff",x"b7",x"6e",x"00",x"00",x"00",x"6e",x"db",x"ff",x"f6",x"ed",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"c4",x"60",x"64",x"b2",x"fb",x"ff",x"ff",x"ff",x"ff",x"fa",x"f1",x"c8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e8",x"e8",x"e8",x"e4",x"e4",x"c4",x"80",x"64",x"d6",x"ff",x"ff",x"92",x"25",x"00",x"01",x"4a",x"db",x"ff",x"fa",x"cd",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"a4",x"80",x"89",x"d6",x"ff",x"ff",x"df",x"ff",x"fb",x"f6",x"ed",x"e8",x"e4",x"e4",x"e8",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e8",x"e4",x"c4",x"80",x"84",x"b2",x"ff",x"ff",x"db",x"49",x"00",x"00",x"00",x"25",x"92",x"fb",x"fb",x"f6",x"cc",x"c4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"a0",x"80",x"84",x"b1",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b2",x"6e",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6e",x"db",x"ff",x"fa",x"f1",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"a0",x"84",x"8d",x"b6",x"fb",x"ff",x"ff",x"ff",x"ff",x"db",x"b7",x"92",x"49",x"00",x"00",x"00",x"00",x"05",x"09",x"0e",x"37",x"5b",x"7b",x"7b",x"5b",x"5b",x"7b",x"7b",x"77",x"97",x"96",x"b2",x"b2",x"ae",x"ad",x"a9",x"a5",x"a5",x"a4",x"a4",x"84",x"80",x"80",x"84",x"a8",x"a9",x"ad",x"ad",x"b2",x"b2",x"b2",x"b6",x"d2",x"d2",x"cd",x"c8",x"c4",x"e4",x"e4",x"c4",x"a4",x"a4",x"f2",x"fb",x"ff",x"72",x"24",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"25",x"49",x"49",x"49",x"6d",x"6d",x"71",x"72",x"72",x"92",x"92",x"96",x"96",x"b6",x"b6",x"b6",x"b6",x"b6",x"ba",x"db",x"db",x"db",x"db",x"db",x"fb",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"20",x"00",x"00",x"00",x"29",x"db",x"ff",x"fa",x"ed",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"ec",x"e8",x"e4",x"e4",x"e8",x"e4",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"84",x"ad",x"d6",x"ff",x"ff",x"b2",x"25",x"00",x"00",x"00",x"45",x"92",x"db",x"ff",x"fa",x"f6",x"ed",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"a4",x"40",x"44",x"b2",x"fb",x"ff",x"ff",x"db",x"73",x"01",x"01",x"49",x"ff",x"fb",x"f1",x"e9",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"a0",x"80",x"a9",x"d6",x"ff",x"ff",x"b7",x"49",x"00",x"01",x"4e",x"bb",x"ff",x"fa",x"f1",x"e8",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"80",x"8d",x"da",x"ff",x"ff",x"ff",x"ff",x"fa",x"f1",x"ed",x"e8",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e8",x"e8",x"e4",x"c4",x"a0",x"80",x"64",x"da",x"ff",x"ff",x"92",x"25",x"00",x"00",x"45",x"b6",x"ff",x"ff",x"f6",x"e9",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"a4",x"64",x"69",x"db",x"ff",x"ff",x"fb",x"ff",x"ff",x"f6",x"ed",x"c4",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"a0",x"84",x"ad",x"fb",x"ff",x"ff",x"49",x"00",x"00",x"49",x"b7",x"ff",x"fa",x"f1",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"c4",x"80",x"84",x"ad",x"fb",x"ff",x"ff",x"ff",x"fb",x"f6",x"f1",x"e9",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"c4",x"a4",x"60",x"89",x"d7",x"ff",x"ff",x"97",x"00",x"00",x"00",x"00",x"4d",x"db",x"fb",x"f6",x"ed",x"c8",x"c4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"c4",x"a4",x"64",x"89",x"db",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"6e",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"96",x"ff",x"fa",x"f1",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"a0",x"80",x"84",x"d6",x"ff",x"ff",x"ff",x"ff",x"ff",x"b7",x"92",x"49",x"00",x"00",x"00",x"00",x"00",x"04",x"09",x"33",x"57",x"5b",x"7b",x"9b",x"9b",x"77",x"77",x"77",x"92",x"6e",x"6d",x"89",x"a9",x"c9",x"c5",x"c5",x"c5",x"c0",x"c0",x"a0",x"80",x"60",x"60",x"64",x"69",x"ae",x"d6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f2",x"c8",x"c4",x"e4",x"e4",x"c4",x"a4",x"ce",x"fb",x"ff",x"92",x"49",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"25",x"6e",x"fb",x"fb",x"f6",x"cd",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"ec",x"e8",x"e4",x"e4",x"e8",x"e4",x"e8",x"e4",x"e4",x"e4",x"e4",x"c4",x"60",x"60",x"d2",x"ff",x"ff",x"d7",x"49",x"00",x"05",x"49",x"92",x"d7",x"fb",x"fb",x"f6",x"f1",x"c8",x"c4",x"c4",x"e4",x"e4",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a4",x"80",x"60",x"69",x"b2",x"fb",x"ff",x"ff",x"db",x"6e",x"05",x"00",x"49",x"b7",x"ff",x"fa",x"ed",x"e8",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"80",x"60",x"b1",x"fb",x"ff",x"db",x"72",x"01",x"00",x"25",x"92",x"df",x"ff",x"f1",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"84",x"b2",x"db",x"ff",x"ff",x"ff",x"ff",x"f6",x"f1",x"e8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e8",x"e8",x"e4",x"e4",x"c4",x"80",x"84",x"8d",x"ff",x"ff",x"fb",x"49",x"00",x"00",x"00",x"6e",x"fb",x"ff",x"fa",x"cd",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e8",x"e4",x"e4",x"e4",x"c4",x"80",x"64",x"91",x"ff",x"ff",x"ff",x"fb",x"ff",x"fa",x"f1",x"c8",x"c4",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"80",x"84",x"d2",x"fb",x"ff",x"bb",x"25",x"00",x"01",x"6e",x"db",x"ff",x"f6",x"f1",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"80",x"a9",x"d6",x"ff",x"df",x"df",x"ff",x"fb",x"f6",x"ed",x"c8",x"c4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"c4",x"a4",x"84",x"b2",x"fb",x"ff",x"bb",x"6e",x"00",x"00",x"00",x"24",x"72",x"ff",x"fb",x"f6",x"ed",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"a0",x"80",x"89",x"b2",x"ff",x"ff",x"df",x"b6",x"6e",x"49",x"25",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"db",x"ff",x"f6",x"ed",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"80",x"84",x"ad",x"fb",x"ff",x"ff",x"db",x"92",x"49",x"25",x"24",x"00",x"00",x"00",x"00",x"04",x"09",x"2d",x"52",x"77",x"77",x"97",x"92",x"b2",x"b2",x"ae",x"8e",x"89",x"a5",x"a5",x"a5",x"c4",x"e5",x"e5",x"e0",x"e4",x"e4",x"c0",x"a0",x"80",x"60",x"64",x"ad",x"b2",x"d6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"cd",x"e4",x"e4",x"e4",x"c4",x"80",x"ad",x"fb",x"ff",x"b6",x"49",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"b7",x"fb",x"fb",x"f1",x"c8",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"60",x"69",x"fb",x"ff",x"ff",x"96",x"49",x"25",x"6e",x"b6",x"fb",x"fb",x"f7",x"f1",x"ed",x"e8",x"c4",x"c4",x"e4",x"e4",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"a0",x"80",x"64",x"48",x"b2",x"fb",x"ff",x"ff",x"db",x"92",x"25",x"00",x"01",x"8e",x"ff",x"ff",x"f6",x"ed",x"c8",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"80",x"84",x"d6",x"ff",x"ff",x"b7",x"49",x"00",x"00",x"49",x"bb",x"ff",x"fa",x"ed",x"c8",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"80",x"84",x"d6",x"ff",x"ff",x"ff",x"ff",x"fb",x"f1",x"ed",x"c8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e8",x"e4",x"c4",x"c4",x"80",x"89",x"d6",x"ff",x"ff",x"b7",x"25",x"00",x"00",x"25",x"92",x"ff",x"fb",x"f5",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"c0",x"80",x"89",x"b6",x"ff",x"ff",x"fb",x"fb",x"fb",x"f6",x"ed",x"c8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"80",x"89",x"d6",x"ff",x"fb",x"92",x"21",x"00",x"25",x"b7",x"fb",x"fb",x"f1",x"cc",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e8",x"e4",x"e4",x"c4",x"a0",x"80",x"d1",x"fb",x"ff",x"df",x"db",x"ff",x"fa",x"f6",x"ed",x"c8",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"84",x"a9",x"d6",x"ff",x"ff",x"96",x"49",x"00",x"00",x"00",x"49",x"b7",x"ff",x"f7",x"f1",x"e8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"60",x"ad",x"fb",x"ff",x"ff",x"b6",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"92",x"ff",x"ff",x"f1",x"cd",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"80",x"84",x"d2",x"fb",x"ff",x"db",x"92",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"4a",x"6e",x"92",x"93",x"92",x"92",x"ae",x"a9",x"a9",x"a9",x"a9",x"c9",x"c4",x"e4",x"e4",x"e0",x"e4",x"e4",x"e0",x"e4",x"c4",x"a0",x"60",x"64",x"89",x"b2",x"d6",x"fb",x"ff",x"ff",x"ff",x"ff",x"df",x"db",x"db",x"bb",x"b7",x"b7",x"ff",x"ff",x"fb",x"ed",x"e8",x"e4",x"e4",x"c0",x"80",x"ad",x"db",x"ff",x"b7",x"49",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"04",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"92",x"fb",x"fb",x"f6",x"cd",x"c8",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e4",x"c4",x"80",x"64",x"b2",x"ff",x"ff",x"df",x"b7",x"96",x"b6",x"db",x"fb",x"fa",x"f2",x"e9",x"e4",x"e4",x"e4",x"e4",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"80",x"60",x"64",x"6d",x"bb",x"db",x"ff",x"ff",x"db",x"92",x"25",x"01",x"01",x"4a",x"b3",x"fb",x"fb",x"f1",x"c8",x"c4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"80",x"64",x"8d",x"fb",x"ff",x"ff",x"6e",x"01",x"00",x"01",x"6e",x"ff",x"ff",x"f6",x"e8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"a0",x"84",x"ad",x"fb",x"ff",x"ff",x"ff",x"ff",x"fb",x"cd",x"c8",x"c4",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"c0",x"a0",x"64",x"ad",x"fb",x"ff",x"db",x"6e",x"00",x"00",x"00",x"4e",x"bb",x"ff",x"fa",x"ed",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"a0",x"60",x"b2",x"fb",x"ff",x"ff",x"fb",x"ff",x"fb",x"f6",x"cc",x"c8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"a0",x"84",x"ad",x"db",x"ff",x"db",x"6e",x"00",x"00",x"4a",x"db",x"ff",x"f6",x"cd",x"c8",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"80",x"84",x"f6",x"ff",x"ff",x"df",x"db",x"fb",x"f6",x"f1",x"c8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"80",x"60",x"d2",x"fb",x"ff",x"db",x"6e",x"00",x"00",x"00",x"00",x"92",x"db",x"ff",x"f6",x"ed",x"e8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"a4",x"60",x"d2",x"fb",x"ff",x"b7",x"6d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"db",x"ff",x"fa",x"cd",x"c8",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"a0",x"80",x"89",x"fa",x"ff",x"ff",x"8e",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"45",x"65",x"ae",x"ae",x"a9",x"89",x"89",x"89",x"84",x"84",x"85",x"cd",x"f2",x"f1",x"ed",x"e9",x"e4",x"e4",x"e0",x"e4",x"c4",x"80",x"40",x"68",x"91",x"d7",x"ff",x"ff",x"ff",x"ff",x"df",x"db",x"b7",x"72",x"4d",x"49",x"49",x"25",x"49",x"b7",x"ff",x"fb",x"cd",x"e8",x"e4",x"e4",x"c0",x"60",x"8d",x"db",x"ff",x"bb",x"4d",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"45",x"45",x"24",x"24",x"24",x"24",x"04",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"b7",x"ff",x"fa",x"f1",x"c8",x"c4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"a0",x"60",x"8d",x"d6",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"f6",x"f2",x"ed",x"e9",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"a4",x"80",x"60",x"60",x"64",x"92",x"bb",x"df",x"ff",x"ff",x"db",x"6e",x"25",x"00",x"00",x"01",x"6e",x"d7",x"ff",x"f6",x"ed",x"c8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"60",x"68",x"b6",x"ff",x"ff",x"db",x"45",x"00",x"00",x"29",x"92",x"ff",x"f6",x"f1",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"80",x"89",x"b6",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"c8",x"c4",x"c4",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"a0",x"80",x"89",x"d6",x"ff",x"ff",x"b7",x"49",x"00",x"00",x"05",x"96",x"df",x"fb",x"f2",x"e8",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"a0",x"80",x"89",x"d6",x"ff",x"ff",x"ff",x"fb",x"ff",x"f6",x"f1",x"c8",x"c4",x"e4",x"e4",x"e8",x"e4",x"e8",x"e8",x"e4",x"e4",x"e4",x"e8",x"e4",x"e4",x"e4",x"c0",x"80",x"89",x"b6",x"ff",x"ff",x"b7",x"45",x"00",x"25",x"92",x"ff",x"fb",x"f1",x"c8",x"c4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"80",x"ad",x"fb",x"ff",x"df",x"df",x"db",x"fb",x"f2",x"cd",x"c4",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"60",x"84",x"d6",x"ff",x"ff",x"b7",x"49",x"00",x"00",x"00",x"25",x"b7",x"fb",x"fb",x"ed",x"e8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"80",x"84",x"d6",x"ff",x"ff",x"92",x"29",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6e",x"ff",x"ff",x"f6",x"c8",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"80",x"84",x"b2",x"ff",x"ff",x"db",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"44",x"69",x"85",x"85",x"84",x"84",x"84",x"60",x"40",x"20",x"40",x"a9",x"f2",x"f6",x"f6",x"f1",x"e8",x"e4",x"e4",x"e4",x"a4",x"60",x"40",x"69",x"b2",x"db",x"ff",x"ff",x"ff",x"df",x"b7",x"72",x"4d",x"29",x"24",x"00",x"00",x"00",x"00",x"05",x"96",x"fb",x"fb",x"cd",x"c4",x"e4",x"e4",x"c0",x"60",x"ad",x"db",x"ff",x"bb",x"6d",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"69",x"69",x"49",x"49",x"49",x"49",x"44",x"24",x"24",x"24",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"6e",x"db",x"ff",x"f6",x"cd",x"c8",x"c4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"c0",x"a0",x"84",x"b2",x"fb",x"ff",x"ff",x"fb",x"fb",x"fa",x"f6",x"ed",x"c8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e8",x"e4",x"e4",x"e4",x"e4",x"c4",x"84",x"64",x"40",x"44",x"69",x"b2",x"db",x"ff",x"ff",x"ff",x"db",x"92",x"25",x"00",x"00",x"00",x"25",x"b2",x"fb",x"fb",x"d1",x"c8",x"e4",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"a0",x"60",x"8d",x"db",x"ff",x"ff",x"b2",x"21",x"00",x"01",x"72",x"db",x"fb",x"f2",x"ed",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"a0",x"60",x"ae",x"db",x"ff",x"ff",x"ff",x"ff",x"f6",x"ed",x"c8",x"c4",x"e4",x"e4",x"e8",x"e8",x"e8",x"e4",x"e8",x"e8",x"e4",x"e4",x"e8",x"e8",x"e4",x"e0",x"e0",x"e4",x"80",x"60",x"b1",x"fb",x"ff",x"db",x"8e",x"01",x"00",x"00",x"29",x"bb",x"ff",x"f6",x"ed",x"e8",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"a0",x"84",x"ad",x"fb",x"ff",x"df",x"ff",x"ff",x"fb",x"f2",x"ec",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"80",x"b2",x"db",x"ff",x"df",x"6e",x"01",x"01",x"4d",x"db",x"ff",x"f6",x"ed",x"c8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"c4",x"80",x"84",x"d2",x"ff",x"ff",x"df",x"df",x"ff",x"fa",x"d1",x"c8",x"c4",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"80",x"80",x"8d",x"db",x"ff",x"df",x"6e",x"04",x"00",x"00",x"00",x"4e",x"db",x"fb",x"f6",x"cd",x"c4",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"60",x"64",x"ad",x"fb",x"ff",x"db",x"6e",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"b6",x"ff",x"fb",x"f1",x"c8",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"a0",x"80",x"89",x"d6",x"ff",x"ff",x"b7",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"24",x"44",x"64",x"40",x"40",x"40",x"40",x"20",x"00",x"00",x"45",x"d2",x"f7",x"f6",x"f2",x"ed",x"c4",x"e4",x"e4",x"c4",x"60",x"40",x"49",x"b6",x"fb",x"ff",x"ff",x"ff",x"bb",x"92",x"4d",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"b6",x"ff",x"fb",x"cd",x"c4",x"e0",x"e0",x"a0",x"80",x"b2",x"ff",x"ff",x"b7",x"49",x"00",x"00",x"00",x"24",x"28",x"49",x"6d",x"6d",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"69",x"69",x"49",x"49",x"49",x"45",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"db",x"ff",x"fb",x"f1",x"c8",x"c4",x"e8",x"e8",x"e8",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"c0",x"a0",x"a8",x"d6",x"ff",x"fa",x"f2",x"f1",x"ed",x"e9",x"e8",x"e4",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"a0",x"80",x"60",x"64",x"6d",x"b6",x"df",x"ff",x"ff",x"ff",x"ff",x"b6",x"69",x"00",x"00",x"00",x"00",x"00",x"49",x"fb",x"fb",x"f6",x"c8",x"c8",x"e8",x"e4",x"e4",x"e4",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"80",x"89",x"b6",x"ff",x"ff",x"d7",x"69",x"00",x"00",x"29",x"b7",x"ff",x"fb",x"ed",x"c8",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"c0",x"a0",x"84",x"b6",x"ff",x"ff",x"ff",x"ff",x"fb",x"f2",x"c8",x"e4",x"e4",x"e4",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"c0",x"80",x"64",x"d6",x"ff",x"ff",x"b6",x"49",x"00",x"00",x"25",x"72",x"df",x"ff",x"f1",x"e8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"a0",x"80",x"89",x"d6",x"ff",x"ff",x"df",x"ff",x"fb",x"f6",x"ed",x"e8",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"80",x"84",x"d6",x"ff",x"ff",x"b7",x"49",x"00",x"29",x"92",x"ff",x"fb",x"f2",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"80",x"80",x"ad",x"fb",x"ff",x"ff",x"db",x"ff",x"ff",x"f6",x"cd",x"c4",x"e4",x"e4",x"e4",x"e4",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"80",x"89",x"d2",x"fb",x"ff",x"db",x"25",x"00",x"00",x"00",x"29",x"96",x"ff",x"fb",x"f1",x"c8",x"c4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"c0",x"60",x"89",x"f7",x"ff",x"ff",x"96",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"92",x"fb",x"fb",x"f6",x"ed",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"80",x"84",x"b2",x"ff",x"ff",x"db",x"6e",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"25",x"6e",x"b7",x"fb",x"f6",x"ed",x"e5",x"c0",x"c0",x"e4",x"c4",x"80",x"40",x"6d",x"bb",x"df",x"ff",x"ff",x"db",x"92",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"d7",x"ff",x"fa",x"c9",x"e4",x"e4",x"e0",x"a0",x"84",x"d6",x"ff",x"ff",x"b6",x"49",x"00",x"00",x"00",x"24",x"49",x"49",x"6d",x"6d",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"72",x"72",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6e",x"ff",x"ff",x"f6",x"ed",x"e8",x"c4",x"e8",x"e8",x"e8",x"e4",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"c0",x"c4",x"cd",x"f6",x"f6",x"f1",x"ed",x"e9",x"c4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"60",x"60",x"64",x"89",x"b2",x"d6",x"ff",x"ff",x"ff",x"ff",x"b7",x"92",x"49",x"00",x"00",x"00",x"00",x"00",x"25",x"92",x"ff",x"fb",x"f1",x"c8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"60",x"ad",x"fb",x"ff",x"df",x"92",x"25",x"00",x"01",x"6e",x"db",x"ff",x"f6",x"c8",x"c4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"80",x"80",x"ad",x"db",x"ff",x"ff",x"ff",x"ff",x"f6",x"ed",x"c4",x"e4",x"e4",x"e4",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"60",x"8d",x"db",x"ff",x"df",x"6e",x"21",x"00",x"00",x"49",x"db",x"ff",x"fa",x"cd",x"e4",x"e4",x"e4",x"e8",x"e8",x"e8",x"e4",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"80",x"84",x"ad",x"fb",x"ff",x"ff",x"df",x"ff",x"fb",x"f2",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"a0",x"80",x"89",x"ff",x"ff",x"df",x"6e",x"01",x"00",x"6e",x"db",x"ff",x"f6",x"ed",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"60",x"84",x"d2",x"ff",x"ff",x"ff",x"db",x"ff",x"fa",x"f1",x"c8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"a4",x"80",x"ad",x"fb",x"ff",x"ff",x"96",x"00",x"00",x"00",x"00",x"6e",x"db",x"ff",x"f6",x"ed",x"c4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"a0",x"64",x"8d",x"fb",x"ff",x"db",x"6e",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"db",x"ff",x"fa",x"f1",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"80",x"89",x"db",x"ff",x"ff",x"92",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"72",x"d7",x"fb",x"f6",x"cd",x"c4",x"e0",x"e0",x"e4",x"c4",x"80",x"60",x"8d",x"d6",x"ff",x"ff",x"df",x"b7",x"6e",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"db",x"fb",x"f6",x"e8",x"e4",x"e4",x"c0",x"a0",x"84",x"d6",x"ff",x"ff",x"92",x"25",x"00",x"00",x"00",x"24",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"96",x"92",x"92",x"72",x"72",x"6d",x"6d",x"4d",x"49",x"49",x"25",x"24",x"24",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"25",x"92",x"ff",x"fa",x"f1",x"e8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e4",x"e4",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"c4",x"ed",x"ed",x"ed",x"e8",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a0",x"80",x"80",x"60",x"40",x"65",x"8d",x"d6",x"fb",x"ff",x"ff",x"ff",x"db",x"b6",x"6d",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"6e",x"d7",x"fb",x"f6",x"ed",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"c0",x"80",x"64",x"d6",x"ff",x"ff",x"b7",x"6a",x"00",x"00",x"25",x"92",x"ff",x"fb",x"f1",x"c8",x"c4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"80",x"84",x"d6",x"ff",x"ff",x"ff",x"ff",x"fb",x"f1",x"e8",x"c4",x"e4",x"e4",x"e4",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"80",x"84",x"b2",x"ff",x"ff",x"bb",x"25",x"00",x"00",x"21",x"92",x"ff",x"fb",x"f1",x"c8",x"e4",x"e4",x"e4",x"e4",x"e8",x"e4",x"e4",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"80",x"88",x"b2",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"ed",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e4",x"c0",x"80",x"84",x"b2",x"ff",x"ff",x"db",x"25",x"00",x"01",x"96",x"ff",x"ff",x"f1",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e4",x"e4",x"80",x"60",x"ad",x"da",x"ff",x"ff",x"ff",x"fb",x"fb",x"f6",x"ed",x"e4",x"e4",x"e8",x"e4",x"e4",x"e4",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a4",x"84",x"88",x"d2",x"ff",x"ff",x"bb",x"6e",x"00",x"00",x"00",x"49",x"b6",x"ff",x"fb",x"f2",x"e8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"80",x"89",x"b6",x"ff",x"ff",x"b7",x"29",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"4e",x"ff",x"ff",x"f6",x"e8",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e4",x"c4",x"80",x"84",x"b2",x"ff",x"ff",x"db",x"6d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"25",x"6e",x"db",x"fb",x"f6",x"cd",x"a4",x"c0",x"e0",x"e4",x"c4",x"60",x"40",x"68",x"da",x"ff",x"ff",x"ff",x"97",x"2d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"6d",x"fb",x"fb",x"f1",x"e4",x"e4",x"e4",x"a0",x"84",x"89",x"fa",x"ff",x"db",x"6d",x"00",x"00",x"00",x"04",x"24",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"96",x"96",x"96",x"92",x"92",x"72",x"6d",x"6d",x"4d",x"49",x"29",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"6e",x"d7",x"fb",x"f6",x"ed",x"e8",x"e4",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e4",x"e9",x"c4",x"c4",x"c0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e4",x"e4",x"e4",x"c4",x"c4",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"60",x"40",x"64",x"89",x"ad",x"b6",x"db",x"fb",x"ff",x"ff",x"ff",x"ff",x"b7",x"6e",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"b2",x"fb",x"fa",x"f1",x"c8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"c0",x"a0",x"60",x"89",x"fb",x"ff",x"ff",x"6e",x"25",x"00",x"01",x"6e",x"db",x"ff",x"f6",x"e9",x"c4",x"c4",x"e8",x"e8",x"e8",x"e4",x"e4",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"a0",x"60",x"89",x"fb",x"ff",x"ff",x"ff",x"ff",x"f6",x"ed",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e4",x"c4",x"a4",x"64",x"ad",x"db",x"ff",x"db",x"92",x"20",x"00",x"00",x"49",x"b7",x"ff",x"f6",x"ed",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"a0",x"84",x"ad",x"db",x"ff",x"ff",x"df",x"ff",x"fa",x"f1",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"a0",x"60",x"8d",x"d6",x"ff",x"ff",x"92",x"00",x"00",x"49",x"db",x"ff",x"f6",x"ed",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"c4",x"80",x"64",x"d6",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"ed",x"c8",x"e4",x"e4",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"80",x"64",x"ad",x"d6",x"ff",x"ff",x"92",x"25",x"00",x"00",x"00",x"92",x"db",x"ff",x"f6",x"ed",x"e8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"c0",x"80",x"64",x"b2",x"db",x"ff",x"db",x"72",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"b7",x"ff",x"fb",x"f1",x"c4",x"e4",x"e8",x"e8",x"e8",x"e4",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"a0",x"80",x"89",x"d6",x"ff",x"ff",x"96",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"b2",x"fb",x"fb",x"f2",x"e9",x"c4",x"e4",x"e4",x"e4",x"a0",x"80",x"40",x"6d",x"b6",x"ff",x"ff",x"fb",x"b2",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"4d",x"b7",x"fb",x"f6",x"ed",x"e4",x"c0",x"c0",x"80",x"84",x"b2",x"ff",x"ff",x"b7",x"49",x"00",x"00",x"00",x"24",x"49",x"49",x"6d",x"6d",x"92",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"24",x"04",x"00",x"00",x"00",x"00",x"00",x"25",x"b3",x"fb",x"fb",x"f1",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"c0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"60",x"64",x"64",x"69",x"6d",x"91",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"4a",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6e",x"db",x"ff",x"f6",x"cd",x"c8",x"e4",x"e4",x"e4",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e4",x"e4",x"a0",x"60",x"64",x"ad",x"ff",x"ff",x"db",x"49",x"00",x"00",x"29",x"92",x"ff",x"fb",x"f2",x"e8",x"e4",x"e4",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"80",x"84",x"b1",x"ff",x"ff",x"ff",x"ff",x"fb",x"f2",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"a0",x"80",x"88",x"b6",x"ff",x"ff",x"b7",x"49",x"00",x"00",x"00",x"92",x"ff",x"ff",x"f2",x"e8",x"e4",x"e4",x"e4",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"80",x"84",x"d6",x"ff",x"ff",x"db",x"db",x"ff",x"fa",x"ed",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"c0",x"a0",x"84",x"b2",x"ff",x"ff",x"d7",x"6a",x"00",x"05",x"72",x"ff",x"ff",x"f6",x"c8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"80",x"89",x"db",x"ff",x"ff",x"df",x"ff",x"ff",x"f2",x"c9",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"60",x"64",x"d6",x"ff",x"ff",x"db",x"49",x"00",x"00",x"00",x"20",x"b7",x"ff",x"fb",x"f1",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"c0",x"80",x"64",x"d6",x"ff",x"ff",x"b7",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6e",x"db",x"fb",x"f6",x"ed",x"e4",x"e4",x"e4",x"e8",x"e4",x"e4",x"e4",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e4",x"c0",x"80",x"84",x"ad",x"fb",x"ff",x"db",x"6e",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"49",x"96",x"fb",x"fb",x"f2",x"e9",x"e4",x"e0",x"e0",x"e4",x"c4",x"80",x"40",x"8d",x"b6",x"ff",x"ff",x"fb",x"d7",x"69",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"72",x"db",x"fb",x"f2",x"e9",x"e0",x"e0",x"a0",x"60",x"64",x"d6",x"ff",x"ff",x"b6",x"25",x"00",x"00",x"00",x"24",x"49",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"d6",x"d6",x"b6",x"b2",x"92",x"8d",x"6d",x"49",x"49",x"44",x"24",x"04",x"00",x"00",x"00",x"00",x"00",x"4a",x"db",x"fb",x"f6",x"ed",x"e8",x"e4",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e4",x"e4",x"e4",x"c4",x"c0",x"e0",x"e0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"c4",x"c4",x"c4",x"c4",x"c0",x"a0",x"80",x"80",x"60",x"60",x"60",x"44",x"48",x"6d",x"92",x"b6",x"db",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b2",x"6e",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"92",x"ff",x"ff",x"d1",x"c8",x"e4",x"e4",x"e4",x"e4",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e4",x"c4",x"a0",x"60",x"89",x"d6",x"ff",x"ff",x"b7",x"01",x"00",x"00",x"6e",x"db",x"ff",x"f6",x"ed",x"e4",x"e4",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"80",x"89",x"d6",x"ff",x"ff",x"ff",x"ff",x"fa",x"f1",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"c0",x"80",x"60",x"ad",x"db",x"ff",x"ff",x"92",x"25",x"00",x"00",x"25",x"db",x"ff",x"f6",x"ed",x"e8",x"e4",x"e4",x"e4",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"80",x"89",x"fb",x"ff",x"ff",x"db",x"db",x"ff",x"f6",x"ed",x"e4",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e4",x"e4",x"e4",x"e0",x"c0",x"a0",x"88",x"d6",x"ff",x"ff",x"b2",x"49",x"00",x"49",x"b7",x"ff",x"fb",x"f1",x"c8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e4",x"e4",x"80",x"84",x"b1",x"ff",x"ff",x"df",x"df",x"ff",x"fb",x"f1",x"c8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"60",x"69",x"fb",x"ff",x"ff",x"92",x"25",x"00",x"00",x"00",x"25",x"db",x"ff",x"f6",x"cd",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"a0",x"84",x"89",x"db",x"ff",x"ff",x"72",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"b6",x"ff",x"fb",x"d1",x"c8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e4",x"a0",x"80",x"89",x"d6",x"ff",x"ff",x"b7",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"4d",x"b6",x"fb",x"fb",x"f2",x"c9",x"e4",x"e0",x"e0",x"e0",x"e0",x"80",x"40",x"64",x"d6",x"ff",x"ff",x"ff",x"d7",x"6e",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"96",x"df",x"f6",x"ed",x"e4",x"e0",x"c0",x"a0",x"60",x"89",x"db",x"ff",x"df",x"92",x"24",x"00",x"00",x"04",x"24",x"49",x"49",x"6d",x"92",x"92",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"6d",x"49",x"49",x"24",x"24",x"04",x"00",x"00",x"00",x"00",x"25",x"b7",x"ff",x"fa",x"f1",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e4",x"c4",x"c0",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"64",x"84",x"85",x"89",x"6d",x"91",x"b2",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b7",x"6e",x"45",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"6e",x"ff",x"fb",x"f6",x"c8",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"c0",x"84",x"64",x"b2",x"ff",x"ff",x"db",x"6e",x"01",x"00",x"01",x"b7",x"ff",x"fb",x"f1",x"e8",x"e4",x"e4",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"a0",x"64",x"b2",x"fb",x"ff",x"ff",x"ff",x"ff",x"f6",x"e9",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"a0",x"60",x"64",x"d6",x"ff",x"ff",x"db",x"49",x"00",x"00",x"25",x"6e",x"db",x"fb",x"f2",x"c8",x"e4",x"e4",x"e4",x"e4",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"60",x"68",x"d6",x"ff",x"ff",x"db",x"ff",x"ff",x"fa",x"f1",x"e4",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e4",x"e4",x"c0",x"a4",x"ad",x"d6",x"ff",x"fb",x"b2",x"6e",x"6e",x"b7",x"ff",x"fb",x"f2",x"e9",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"a4",x"60",x"89",x"fb",x"ff",x"ff",x"bf",x"ff",x"fb",x"f1",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"80",x"89",x"b2",x"ff",x"ff",x"d7",x"49",x"01",x"00",x"00",x"25",x"92",x"ff",x"fb",x"f1",x"c8",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"60",x"84",x"d2",x"ff",x"ff",x"db",x"29",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"92",x"db",x"ff",x"f6",x"cd",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"c0",x"c4",x"80",x"60",x"b2",x"fb",x"ff",x"db",x"72",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"8e",x"db",x"fb",x"f6",x"cd",x"c8",x"e4",x"e0",x"e0",x"e4",x"c4",x"a0",x"40",x"68",x"b2",x"fb",x"ff",x"ff",x"b7",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"b6",x"fb",x"fa",x"c9",x"e4",x"e4",x"e4",x"a0",x"60",x"89",x"b2",x"fb",x"ff",x"bb",x"25",x"00",x"00",x"00",x"24",x"25",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"4a",x"db",x"ff",x"f6",x"ec",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"c0",x"a0",x"a0",x"84",x"60",x"64",x"64",x"84",x"84",x"84",x"64",x"64",x"64",x"69",x"89",x"8d",x"8d",x"b2",x"b2",x"b6",x"ba",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b7",x"96",x"6e",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"29",x"92",x"ff",x"fb",x"f1",x"c4",x"e4",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e4",x"e4",x"a0",x"60",x"89",x"d6",x"ff",x"ff",x"b7",x"29",x"00",x"01",x"49",x"db",x"ff",x"f6",x"ed",x"e4",x"e4",x"e4",x"e4",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"c0",x"80",x"69",x"d6",x"ff",x"ff",x"ff",x"ff",x"fa",x"f1",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"c0",x"80",x"84",x"8d",x"fb",x"ff",x"ff",x"92",x"25",x"00",x"00",x"49",x"b7",x"ff",x"fb",x"ed",x"c4",x"c4",x"e4",x"e4",x"e4",x"e4",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"64",x"8d",x"fb",x"ff",x"ff",x"db",x"ff",x"fb",x"f2",x"e9",x"e4",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e4",x"e4",x"e0",x"c0",x"c4",x"cd",x"f6",x"fb",x"fb",x"d7",x"b6",x"d7",x"fb",x"ff",x"f6",x"ed",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"64",x"b1",x"ff",x"ff",x"df",x"bf",x"ff",x"fa",x"ed",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"a0",x"80",x"ad",x"db",x"ff",x"fb",x"b2",x"21",x"00",x"00",x"00",x"4d",x"d7",x"ff",x"f6",x"ed",x"c4",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e4",x"c4",x"a0",x"60",x"ad",x"fb",x"ff",x"df",x"b6",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"d7",x"ff",x"fa",x"f1",x"c8",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"80",x"84",x"d6",x"ff",x"ff",x"b7",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"8e",x"d7",x"fb",x"f6",x"f1",x"c4",x"c0",x"e0",x"e0",x"e4",x"c4",x"a0",x"60",x"44",x"91",x"fb",x"ff",x"ff",x"db",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"6e",x"fb",x"fb",x"f1",x"c4",x"e0",x"e4",x"c4",x"80",x"40",x"ad",x"db",x"ff",x"ff",x"96",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"6d",x"6d",x"92",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"25",x"92",x"fb",x"fb",x"f1",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"80",x"a9",x"ad",x"ad",x"ad",x"b2",x"b2",x"b2",x"b2",x"d6",x"d6",x"d6",x"db",x"db",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"6d",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"d7",x"fb",x"f6",x"ed",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e4",x"e4",x"80",x"60",x"b1",x"fb",x"ff",x"db",x"6e",x"00",x"00",x"25",x"92",x"fb",x"fb",x"f2",x"e9",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"a0",x"84",x"8d",x"db",x"ff",x"ff",x"ff",x"ff",x"f6",x"ed",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"c0",x"80",x"a8",x"d2",x"ff",x"ff",x"db",x"69",x"20",x"00",x"00",x"6e",x"db",x"ff",x"f6",x"ed",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e4",x"c0",x"80",x"89",x"b2",x"fb",x"ff",x"ff",x"ff",x"ff",x"fb",x"cd",x"c4",x"c4",x"e4",x"e4",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"c4",x"e4",x"e9",x"f1",x"f6",x"fb",x"fb",x"fb",x"f7",x"fb",x"f6",x"ed",x"e8",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e4",x"a0",x"60",x"a9",x"d6",x"ff",x"fb",x"df",x"df",x"fb",x"f6",x"ed",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"a0",x"80",x"84",x"b2",x"ff",x"ff",x"db",x"6e",x"00",x"00",x"00",x"25",x"92",x"fb",x"fb",x"f6",x"e8",x"c4",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"80",x"88",x"d2",x"ff",x"ff",x"d7",x"6d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"49",x"92",x"ff",x"fb",x"f6",x"c9",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e4",x"e4",x"80",x"84",x"ad",x"fb",x"ff",x"ff",x"92",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"92",x"db",x"fb",x"f6",x"cd",x"c8",x"c0",x"c0",x"e0",x"e4",x"c4",x"a4",x"60",x"60",x"8d",x"db",x"ff",x"ff",x"db",x"92",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"69",x"d7",x"ff",x"f6",x"c9",x"e4",x"e4",x"e0",x"a0",x"80",x"64",x"b2",x"fb",x"ff",x"db",x"6e",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"6d",x"6d",x"49",x"49",x"24",x"20",x"00",x"00",x"00",x"00",x"6e",x"db",x"fb",x"f6",x"ed",x"c8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e4",x"e4",x"a0",x"80",x"89",x"d6",x"fb",x"fb",x"fb",x"fb",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b7",x"92",x"6d",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"b2",x"fb",x"f7",x"f2",x"e9",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"a4",x"60",x"64",x"fb",x"ff",x"fb",x"8e",x"25",x"00",x"00",x"6d",x"db",x"fb",x"f6",x"cd",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e4",x"e4",x"e0",x"e0",x"e4",x"e4",x"e0",x"c0",x"80",x"84",x"b6",x"ff",x"ff",x"ff",x"ff",x"fb",x"f1",x"c8",x"c0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"60",x"ad",x"fb",x"ff",x"ff",x"92",x"00",x"00",x"00",x"49",x"b6",x"ff",x"fb",x"f2",x"c8",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e4",x"a0",x"80",x"ad",x"db",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"c9",x"c4",x"e0",x"e4",x"e4",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e9",x"e9",x"ed",x"ee",x"ee",x"ed",x"e9",x"e9",x"e4",x"c4",x"c0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"80",x"60",x"d2",x"fb",x"ff",x"ff",x"ff",x"ff",x"f6",x"f1",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"c0",x"80",x"80",x"a9",x"db",x"ff",x"ff",x"92",x"25",x"00",x"00",x"25",x"92",x"d7",x"fb",x"f6",x"ed",x"e4",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"80",x"ad",x"db",x"ff",x"ff",x"92",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"49",x"92",x"db",x"fb",x"fb",x"f2",x"c9",x"c4",x"c0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"c0",x"60",x"84",x"d2",x"ff",x"ff",x"b7",x"29",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"8e",x"b6",x"fb",x"fb",x"f6",x"cd",x"c4",x"c0",x"e0",x"e0",x"e0",x"c4",x"a0",x"40",x"64",x"8d",x"d7",x"ff",x"ff",x"ff",x"92",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"b6",x"fb",x"f6",x"cd",x"c4",x"e4",x"e4",x"c0",x"80",x"84",x"8d",x"db",x"ff",x"ff",x"92",x"25",x"00",x"00",x"00",x"00",x"24",x"49",x"6d",x"6d",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"6d",x"6d",x"49",x"28",x"24",x"20",x"00",x"00",x"00",x"04",x"96",x"ff",x"fb",x"f1",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e4",x"c0",x"80",x"88",x"b2",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"db",x"db",x"db",x"bb",x"b7",x"b6",x"92",x"92",x"6e",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"d7",x"fb",x"f2",x"ed",x"c4",x"e4",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"c0",x"80",x"64",x"8d",x"ff",x"ff",x"db",x"69",x"25",x"24",x"49",x"b6",x"ff",x"f7",x"f2",x"c8",x"c4",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"e4",x"c0",x"80",x"60",x"8d",x"db",x"ff",x"ff",x"ff",x"ff",x"f6",x"c9",x"c4",x"c0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"a0",x"84",x"b1",x"ff",x"ff",x"bb",x"6e",x"00",x"24",x"49",x"92",x"db",x"fb",x"f2",x"cd",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"c0",x"80",x"64",x"d2",x"ff",x"ff",x"ff",x"ff",x"ff",x"f6",x"ed",x"c4",x"c0",x"e0",x"e4",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e4",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e9",x"c4",x"c4",x"c4",x"e0",x"e4",x"e4",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"a0",x"80",x"88",x"fb",x"ff",x"ff",x"ff",x"ff",x"fb",x"f2",x"e9",x"e4",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"c0",x"80",x"84",x"d1",x"ff",x"ff",x"df",x"4e",x"04",x"25",x"29",x"6d",x"db",x"fb",x"f6",x"ed",x"e8",x"e4",x"c0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"c0",x"a0",x"84",x"d6",x"ff",x"ff",x"bb",x"6d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"45",x"6e",x"b2",x"fb",x"fb",x"f6",x"f1",x"c9",x"c4",x"c0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"c0",x"80",x"a9",x"fb",x"ff",x"df",x"72",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"25",x"49",x"b2",x"d7",x"fb",x"f7",x"f2",x"e9",x"c4",x"c0",x"e0",x"e0",x"e0",x"c0",x"a0",x"60",x"44",x"8d",x"d6",x"ff",x"ff",x"ff",x"b2",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"29",x"b6",x"fb",x"fa",x"cd",x"c4",x"c0",x"e4",x"c0",x"a0",x"80",x"89",x"d6",x"ff",x"ff",x"db",x"49",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"6d",x"91",x"92",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"24",x"24",x"20",x"00",x"00",x"00",x"29",x"db",x"ff",x"f6",x"e9",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e4",x"a0",x"60",x"ad",x"db",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"b7",x"b6",x"92",x"92",x"6e",x"6d",x"69",x"49",x"25",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"92",x"fb",x"fb",x"ed",x"c4",x"c4",x"e0",x"e0",x"e4",x"e0",x"e0",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"88",x"b6",x"ff",x"ff",x"db",x"6d",x"49",x"72",x"b6",x"fb",x"fb",x"f2",x"e9",x"c4",x"c0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"60",x"64",x"b2",x"ff",x"ff",x"ff",x"ff",x"fb",x"f1",x"c4",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"a4",x"a8",x"d6",x"ff",x"df",x"97",x"4e",x"49",x"6e",x"d6",x"fb",x"fb",x"f2",x"cd",x"c4",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e4",x"e0",x"e0",x"c0",x"a0",x"84",x"89",x"db",x"ff",x"ff",x"df",x"df",x"fb",x"f2",x"e9",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e4",x"c0",x"80",x"84",x"ad",x"ff",x"ff",x"df",x"ff",x"ff",x"fa",x"ed",x"c8",x"e4",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"c0",x"80",x"a8",x"f6",x"ff",x"df",x"b7",x"4d",x"49",x"92",x"b6",x"db",x"fb",x"f6",x"ed",x"c4",x"c4",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"c0",x"a0",x"84",x"fa",x"ff",x"df",x"92",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"8e",x"b7",x"f7",x"fb",x"fb",x"f2",x"cd",x"c4",x"c0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"a0",x"a4",x"d2",x"ff",x"ff",x"bb",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"29",x"6d",x"92",x"d6",x"fb",x"fb",x"f2",x"c9",x"c4",x"c4",x"c0",x"e0",x"e0",x"e0",x"e4",x"a0",x"60",x"44",x"8d",x"b6",x"ff",x"ff",x"ff",x"b7",x"29",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"92",x"fb",x"fb",x"f2",x"c4",x"c0",x"e4",x"e0",x"a0",x"80",x"84",x"ae",x"fb",x"ff",x"df",x"92",x"24",x"00",x"00",x"00",x"00",x"24",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"92",x"6d",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"05",x"72",x"ff",x"ff",x"f2",x"e8",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e4",x"e4",x"e4",x"c0",x"80",x"80",x"d2",x"ff",x"df",x"bb",x"92",x"6e",x"49",x"45",x"45",x"45",x"25",x"25",x"25",x"25",x"24",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"d7",x"fb",x"f6",x"c9",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"cd",x"f6",x"ff",x"ff",x"ff",x"b6",x"b6",x"d6",x"fb",x"f6",x"f2",x"e9",x"e4",x"e4",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"60",x"8d",x"db",x"ff",x"ff",x"ff",x"ff",x"f6",x"e9",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"c0",x"c4",x"cd",x"fa",x"ff",x"df",x"bb",x"b7",x"d7",x"d7",x"f7",x"f6",x"f2",x"e9",x"c4",x"c4",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e4",x"e0",x"e0",x"c0",x"80",x"84",x"b2",x"ff",x"ff",x"df",x"df",x"fb",x"fa",x"ed",x"e4",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e4",x"e4",x"a0",x"60",x"89",x"d6",x"ff",x"ff",x"db",x"ff",x"fb",x"f2",x"e9",x"c4",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"c4",x"a0",x"c9",x"f6",x"ff",x"ff",x"db",x"d6",x"d6",x"fb",x"fb",x"f6",x"f2",x"c9",x"e4",x"e4",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"c0",x"a4",x"a9",x"fb",x"ff",x"df",x"4d",x"00",x"00",x"00",x"00",x"25",x"69",x"8e",x"b2",x"d6",x"f7",x"f6",x"f6",x"f2",x"cd",x"c4",x"c0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"c0",x"a0",x"c9",x"f6",x"ff",x"df",x"92",x"05",x"00",x"00",x"01",x"25",x"49",x"6d",x"92",x"b6",x"d7",x"f7",x"f6",x"f2",x"e9",x"e5",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"60",x"64",x"8d",x"d7",x"ff",x"ff",x"ff",x"b7",x"6d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"92",x"d7",x"f6",x"f2",x"e9",x"c0",x"e0",x"e4",x"c0",x"80",x"60",x"ad",x"d6",x"ff",x"ff",x"b7",x"49",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"6d",x"91",x"92",x"92",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"49",x"b7",x"ff",x"fa",x"ed",x"e4",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e4",x"e4",x"e4",x"a0",x"80",x"89",x"db",x"ff",x"df",x"72",x"29",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"72",x"fb",x"f7",x"ee",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"e9",x"f6",x"fb",x"ff",x"fb",x"f6",x"f6",x"f6",x"f2",x"ed",x"e9",x"e4",x"e0",x"e4",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"e4",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"64",x"b2",x"ff",x"ff",x"ff",x"ff",x"fb",x"ed",x"e4",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e4",x"ed",x"f6",x"fb",x"ff",x"fb",x"fb",x"f7",x"f2",x"f2",x"ed",x"e9",x"e4",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"89",x"d6",x"ff",x"ff",x"db",x"ff",x"fb",x"f6",x"e9",x"c0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e4",x"c4",x"a0",x"60",x"8d",x"db",x"df",x"df",x"df",x"ff",x"fb",x"ed",x"c4",x"c0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e4",x"c4",x"c8",x"f6",x"fb",x"fb",x"f7",x"fb",x"fb",x"f6",x"f2",x"ed",x"c8",x"c4",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"c0",x"c4",x"c9",x"fa",x"ff",x"db",x"6e",x"49",x"49",x"49",x"6d",x"8e",x"b2",x"f6",x"fb",x"f6",x"f6",x"f2",x"ed",x"c9",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"c4",x"c9",x"f6",x"ff",x"ff",x"96",x"49",x"49",x"4a",x"6e",x"8e",x"b2",x"d6",x"f7",x"fb",x"f6",x"f2",x"ed",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"a0",x"60",x"40",x"8d",x"b6",x"ff",x"ff",x"ff",x"db",x"6e",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"92",x"db",x"fb",x"f2",x"e9",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"64",x"d6",x"ff",x"ff",x"db",x"72",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"04",x"92",x"fb",x"fb",x"f2",x"e8",x"e4",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"80",x"84",x"d2",x"ff",x"ff",x"df",x"4d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"b6",x"ff",x"f6",x"e9",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"ed",x"f2",x"f6",x"f2",x"f2",x"ed",x"e9",x"e4",x"e4",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"80",x"60",x"89",x"db",x"ff",x"ff",x"ff",x"ff",x"f6",x"e9",x"e4",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"ed",x"f2",x"f2",x"f6",x"f2",x"ed",x"e9",x"e4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"ad",x"ff",x"ff",x"ff",x"fb",x"fb",x"fa",x"f1",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"89",x"d2",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"e9",x"c4",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e4",x"e4",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e4",x"c0",x"c4",x"ed",x"f2",x"f6",x"f2",x"f2",x"ed",x"c9",x"c4",x"c4",x"c4",x"e4",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c4",x"e9",x"f2",x"fa",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"f6",x"f6",x"f2",x"ed",x"ed",x"c9",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"c4",x"c8",x"f1",x"fa",x"ff",x"ff",x"d7",x"d7",x"d7",x"fb",x"fb",x"fb",x"f7",x"f2",x"f2",x"c9",x"e5",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"c4",x"a4",x"40",x"40",x"8d",x"d6",x"ff",x"ff",x"ff",x"d7",x"6e",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"92",x"fb",x"fb",x"f6",x"e9",x"c0",x"c0",x"e0",x"c0",x"a0",x"80",x"84",x"ad",x"fb",x"ff",x"ff",x"96",x"29",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"49",x"b7",x"fb",x"f6",x"ed",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"89",x"fb",x"ff",x"ff",x"b7",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6e",x"db",x"fb",x"f2",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c4",x"c8",x"c8",x"c4",x"e4",x"e0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"60",x"64",x"b2",x"fb",x"ff",x"ff",x"ff",x"fb",x"f2",x"e4",x"e0",x"e0",x"e0",x"e0",x"e4",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e8",x"e9",x"c4",x"c4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a4",x"d2",x"ff",x"ff",x"ff",x"fb",x"fa",x"f2",x"e8",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"c0",x"a0",x"a0",x"c0",x"e0",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"a0",x"ad",x"f6",x"ff",x"ff",x"ff",x"ff",x"f6",x"ed",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e4",x"e8",x"e9",x"c9",x"e9",x"e4",x"e4",x"e4",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"ed",x"f2",x"f6",x"f6",x"f6",x"f6",x"f6",x"f2",x"f2",x"ed",x"ed",x"c8",x"c4",x"c4",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"c4",x"c9",x"f1",x"f6",x"f6",x"f6",x"f2",x"f2",x"f2",x"f2",x"ee",x"c9",x"c9",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e4",x"e0",x"e0",x"e4",x"c4",x"80",x"60",x"64",x"8d",x"da",x"ff",x"ff",x"ff",x"b7",x"69",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"b2",x"fb",x"fb",x"f2",x"e9",x"e4",x"c0",x"c0",x"e0",x"a0",x"60",x"64",x"8d",x"da",x"ff",x"ff",x"db",x"49",x"00",x"00",x"00",x"00",x"04",x"24",x"49",x"49",x"6d",x"6d",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"92",x"fb",x"fb",x"f2",x"c8",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"88",x"b2",x"ff",x"ff",x"db",x"6e",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"92",x"fb",x"fb",x"cd",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"60",x"8d",x"d6",x"ff",x"ff",x"fb",x"ff",x"fb",x"cd",x"c4",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e0",x"e0",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"c9",x"f6",x"ff",x"ff",x"ff",x"fb",x"f6",x"ed",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"a0",x"80",x"80",x"a4",x"a4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"d2",x"fb",x"ff",x"ff",x"ff",x"fb",x"f2",x"e9",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e4",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e4",x"e8",x"e9",x"e9",x"ed",x"ed",x"e9",x"e9",x"e9",x"e8",x"e4",x"c4",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"e0",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c4",x"e8",x"e9",x"ed",x"ed",x"e9",x"e9",x"e9",x"e9",x"e4",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e0",x"c0",x"a0",x"80",x"60",x"44",x"91",x"db",x"ff",x"ff",x"ff",x"d7",x"69",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"92",x"fb",x"fb",x"f2",x"e9",x"e0",x"e0",x"e0",x"c0",x"c0",x"80",x"60",x"89",x"b6",x"ff",x"ff",x"db",x"92",x"25",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"6d",x"6d",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"04",x"d7",x"ff",x"f7",x"c9",x"c4",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"a0",x"60",x"ad",x"da",x"ff",x"ff",x"b7",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"b7",x"fb",x"f6",x"c9",x"c4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"64",x"91",x"ff",x"ff",x"fb",x"fb",x"fb",x"f6",x"c9",x"c0",x"e0",x"e0",x"e0",x"e4",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"c0",x"a0",x"ee",x"fb",x"ff",x"ff",x"ff",x"fa",x"ed",x"c4",x"c0",x"e0",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"60",x"88",x"ad",x"a9",x"a4",x"a0",x"a0",x"a0",x"a0",x"c0",x"a0",x"a0",x"80",x"60",x"60",x"80",x"80",x"a4",x"c4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e0",x"e0",x"e0",x"c0",x"a0",x"ce",x"fb",x"ff",x"ff",x"fb",x"f2",x"c9",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"c0",x"c0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c4",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"a0",x"60",x"60",x"68",x"b2",x"db",x"ff",x"ff",x"ff",x"b7",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"69",x"b7",x"fb",x"f7",x"d2",x"c9",x"e0",x"e0",x"e0",x"e0",x"c4",x"80",x"60",x"64",x"b6",x"df",x"ff",x"ff",x"b2",x"45",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"6d",x"6d",x"92",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"92",x"92",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"24",x"6d",x"fb",x"fb",x"f2",x"c8",x"c4",x"c0",x"e0",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"60",x"b2",x"ff",x"ff",x"db",x"6e",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"b6",x"fb",x"f2",x"a4",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"60",x"89",x"d6",x"ff",x"fb",x"fb",x"ff",x"fb",x"f2",x"c9",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e0",x"c0",x"c4",x"ed",x"f6",x"fb",x"fa",x"f6",x"f1",x"c8",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"c0",x"a0",x"60",x"64",x"8d",x"b6",x"d6",x"d2",x"ad",x"84",x"80",x"60",x"60",x"60",x"60",x"60",x"64",x"64",x"69",x"ad",x"cd",x"c9",x"c4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a4",x"ed",x"f6",x"fb",x"f6",x"f2",x"e9",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e0",x"c0",x"a0",x"a0",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"80",x"60",x"80",x"a0",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"c0",x"c0",x"a0",x"80",x"60",x"60",x"89",x"b2",x"db",x"ff",x"ff",x"df",x"b6",x"4d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"4e",x"b6",x"fb",x"f6",x"ed",x"e9",x"e4",x"e0",x"e0",x"e0",x"c0",x"80",x"40",x"64",x"b2",x"db",x"ff",x"ff",x"b6",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"48",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"da",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"6d",x"6d",x"49",x"28",x"24",x"00",x"00",x"00",x"00",x"49",x"b7",x"fb",x"f6",x"ed",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"a0",x"80",x"68",x"b6",x"ff",x"ff",x"b2",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"24",x"24",x"24",x"25",x"25",x"25",x"25",x"25",x"25",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"fb",x"d2",x"89",x"60",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"60",x"b2",x"fb",x"ff",x"d7",x"db",x"ff",x"fb",x"ee",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c4",x"c8",x"ed",x"f2",x"f1",x"ed",x"e8",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a4",x"80",x"60",x"64",x"8d",x"b6",x"ff",x"ff",x"db",x"b6",x"8d",x"8d",x"69",x"69",x"69",x"69",x"69",x"8d",x"92",x"b6",x"d6",x"f6",x"f2",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c4",x"e9",x"ed",x"f1",x"ed",x"e9",x"e4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"84",x"c4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"40",x"64",x"a9",x"c9",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"40",x"64",x"8d",x"d6",x"fb",x"ff",x"ff",x"db",x"96",x"49",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"6e",x"b7",x"fb",x"f6",x"cd",x"c4",x"e4",x"e0",x"e0",x"e0",x"c0",x"80",x"60",x"64",x"92",x"db",x"ff",x"ff",x"db",x"6d",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"6e",x"d7",x"fb",x"f2",x"e9",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"84",x"b1",x"db",x"ff",x"db",x"6e",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"25",x"29",x"49",x"6d",x"8e",x"8e",x"8e",x"92",x"b2",x"b2",x"d6",x"d7",x"d7",x"d7",x"f7",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"ff",x"ff",x"fb",x"b2",x"8d",x"ad",x"ad",x"a9",x"a9",x"a9",x"89",x"88",x"84",x"84",x"84",x"84",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"80",x"64",x"d6",x"ff",x"ff",x"96",x"96",x"df",x"fb",x"f2",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"80",x"a4",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e9",x"e4",x"c4",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"84",x"ad",x"da",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"d7",x"f7",x"f7",x"fb",x"fb",x"db",x"ff",x"ff",x"ff",x"fb",x"d2",x"a4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c4",x"c4",x"c4",x"c0",x"c0",x"e0",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"60",x"60",x"64",x"89",x"ad",x"d1",x"cd",x"c4",x"c0",x"c0",x"e0",x"e4",x"e4",x"e4",x"e0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"80",x"60",x"60",x"89",x"d2",x"fb",x"f6",x"f2",x"c4",x"c0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"c0",x"80",x"60",x"60",x"69",x"8e",x"d6",x"fb",x"ff",x"ff",x"ff",x"db",x"72",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"b2",x"fb",x"fb",x"f6",x"c9",x"a4",x"c0",x"e0",x"e0",x"e0",x"c0",x"a0",x"60",x"64",x"d2",x"fb",x"ff",x"ff",x"db",x"6e",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"92",x"92",x"92",x"6d",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"45",x"b2",x"fb",x"f6",x"ed",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"89",x"d6",x"ff",x"ff",x"b7",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"45",x"49",x"69",x"6d",x"6e",x"92",x"92",x"b6",x"b7",x"db",x"db",x"db",x"db",x"db",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"f7",x"fb",x"fb",x"fb",x"fb",x"d6",x"d2",x"d2",x"d2",x"d2",x"d2",x"d2",x"d2",x"d2",x"b2",x"b1",x"b1",x"ad",x"ad",x"ad",x"a9",x"a9",x"a9",x"a9",x"a4",x"a4",x"a4",x"84",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"80",x"89",x"fb",x"ff",x"db",x"6e",x"72",x"df",x"fb",x"f2",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"64",x"69",x"ad",x"cd",x"c9",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"c4",x"a0",x"80",x"60",x"60",x"88",x"ad",x"d6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"d6",x"a9",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"60",x"69",x"ad",x"d6",x"fa",x"fb",x"d2",x"c9",x"a4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"60",x"60",x"64",x"89",x"b2",x"fb",x"ff",x"ff",x"f6",x"c9",x"a4",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"64",x"69",x"92",x"db",x"ff",x"ff",x"ff",x"ff",x"d7",x"6e",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"6d",x"b6",x"f7",x"f6",x"f2",x"e9",x"c4",x"c0",x"c0",x"e0",x"e4",x"c0",x"a0",x"60",x"64",x"ad",x"fb",x"ff",x"ff",x"db",x"72",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"48",x"49",x"6d",x"6d",x"6d",x"92",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"6e",x"d7",x"fb",x"f2",x"c9",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"60",x"ad",x"fb",x"ff",x"db",x"92",x"25",x"00",x"01",x"01",x"01",x"21",x"49",x"6e",x"8e",x"92",x"b6",x"d7",x"db",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"f6",x"f6",x"f6",x"f6",x"f2",x"f2",x"f1",x"f1",x"ed",x"ed",x"ed",x"ed",x"ed",x"ed",x"ed",x"ed",x"ed",x"ed",x"ed",x"ed",x"ee",x"ee",x"ed",x"ed",x"f2",x"f2",x"f2",x"f2",x"f2",x"f6",x"f6",x"f6",x"f6",x"f6",x"f6",x"f6",x"f6",x"f6",x"f2",x"f2",x"f2",x"d2",x"cd",x"cd",x"ad",x"a9",x"89",x"84",x"64",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"84",x"d2",x"ff",x"df",x"92",x"25",x"4d",x"df",x"ff",x"f6",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"80",x"60",x"40",x"64",x"8d",x"b6",x"db",x"fb",x"f2",x"c9",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a4",x"a0",x"80",x"60",x"64",x"89",x"b2",x"fb",x"ff",x"ff",x"ff",x"bb",x"b7",x"b7",x"db",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"df",x"ff",x"ff",x"fb",x"ce",x"c4",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"60",x"64",x"8d",x"b6",x"db",x"ff",x"ff",x"ff",x"fa",x"cd",x"a9",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"60",x"60",x"69",x"92",x"d6",x"fb",x"ff",x"ff",x"ff",x"fb",x"d2",x"a9",x"a4",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c4",x"c0",x"a0",x"80",x"60",x"60",x"64",x"8d",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"b7",x"6e",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"6e",x"d7",x"fb",x"f6",x"ed",x"e8",x"c0",x"e0",x"e0",x"e0",x"c0",x"c4",x"a0",x"60",x"60",x"8d",x"db",x"ff",x"ff",x"ff",x"92",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"8d",x"6d",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"b6",x"fb",x"f7",x"ed",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"89",x"b6",x"ff",x"ff",x"bb",x"92",x"49",x"49",x"8e",x"b2",x"b7",x"d7",x"fb",x"fb",x"fb",x"fb",x"fb",x"f7",x"f7",x"f6",x"f2",x"f2",x"f2",x"ee",x"ed",x"e9",x"e9",x"e9",x"e9",x"e5",x"c4",x"c4",x"c4",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"c0",x"c0",x"c4",x"c4",x"c4",x"c4",x"c9",x"c9",x"c9",x"ed",x"ed",x"ed",x"f2",x"f2",x"f2",x"f2",x"f2",x"f2",x"f6",x"f6",x"f6",x"f6",x"f6",x"f6",x"f6",x"d2",x"d2",x"b1",x"ad",x"ad",x"ad",x"a9",x"88",x"84",x"84",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"a0",x"60",x"ad",x"fb",x"ff",x"b7",x"49",x"00",x"49",x"df",x"ff",x"f6",x"c9",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"60",x"60",x"64",x"69",x"b2",x"da",x"fb",x"ff",x"ff",x"ff",x"fb",x"ce",x"a4",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"60",x"60",x"64",x"8d",x"d6",x"db",x"ff",x"ff",x"ff",x"db",x"92",x"49",x"25",x"00",x"05",x"49",x"6e",x"92",x"92",x"92",x"6e",x"72",x"6e",x"29",x"4d",x"b6",x"ff",x"ff",x"f6",x"c9",x"a0",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a0",x"60",x"40",x"64",x"89",x"ad",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d2",x"a9",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"60",x"40",x"64",x"8d",x"d6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"f6",x"cd",x"80",x"a0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"60",x"60",x"60",x"64",x"89",x"b2",x"d6",x"fb",x"ff",x"ff",x"ff",x"ff",x"b7",x"6e",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"6e",x"d7",x"fb",x"f7",x"f2",x"c9",x"c4",x"c0",x"e0",x"e0",x"e0",x"e4",x"c4",x"80",x"60",x"64",x"b2",x"db",x"ff",x"ff",x"db",x"92",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"6d",x"49",x"49",x"29",x"24",x"00",x"00",x"00",x"00",x"49",x"db",x"fb",x"f2",x"c9",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"b1",x"db",x"ff",x"ff",x"db",x"b6",x"b2",x"b2",x"d7",x"f7",x"fb",x"fb",x"fb",x"f6",x"f6",x"f2",x"f2",x"ee",x"ed",x"e9",x"e9",x"e9",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e9",x"e9",x"e9",x"e9",x"ed",x"ed",x"f1",x"f2",x"f2",x"f2",x"f6",x"f6",x"f6",x"f6",x"f6",x"d6",x"d6",x"d6",x"d6",x"d2",x"d1",x"ad",x"ad",x"a9",x"a9",x"a4",x"84",x"84",x"84",x"a0",x"a0",x"80",x"80",x"60",x"64",x"b2",x"ff",x"db",x"6e",x"01",x"00",x"25",x"b7",x"ff",x"fb",x"f2",x"c9",x"a0",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"84",x"89",x"8d",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"f6",x"cd",x"a4",x"a0",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"60",x"64",x"8d",x"b2",x"da",x"ff",x"ff",x"ff",x"ff",x"db",x"6e",x"29",x"00",x"00",x"00",x"00",x"00",x"25",x"25",x"25",x"25",x"25",x"25",x"24",x"00",x"04",x"4d",x"db",x"ff",x"fb",x"d2",x"a9",x"a4",x"a0",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"80",x"a4",x"c4",x"c4",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"64",x"6d",x"b2",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"db",x"b7",x"db",x"ff",x"ff",x"fb",x"d2",x"a9",x"a0",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a0",x"80",x"80",x"60",x"64",x"89",x"8d",x"b2",x"db",x"ff",x"ff",x"ff",x"ff",x"fb",x"d7",x"92",x"b7",x"df",x"ff",x"ff",x"f6",x"a9",x"a0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"60",x"44",x"64",x"89",x"b2",x"b6",x"fb",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"92",x"db",x"fb",x"f7",x"ee",x"c5",x"c0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"80",x"60",x"64",x"b1",x"fb",x"ff",x"ff",x"df",x"92",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"49",x"49",x"24",x"04",x"00",x"00",x"00",x"25",x"92",x"ff",x"f7",x"cd",x"a4",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"80",x"d6",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"f7",x"f6",x"f6",x"f2",x"f2",x"ed",x"e9",x"c9",x"c9",x"c4",x"c4",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c4",x"c4",x"c4",x"e8",x"e9",x"e9",x"ed",x"ed",x"f1",x"f2",x"f6",x"f6",x"f6",x"f6",x"f6",x"f6",x"f6",x"f6",x"f6",x"f6",x"d2",x"cd",x"ad",x"a9",x"84",x"84",x"60",x"40",x"40",x"89",x"d6",x"ff",x"b7",x"4a",x"01",x"00",x"25",x"6e",x"db",x"ff",x"fb",x"d2",x"a9",x"80",x"80",x"a0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"89",x"8d",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"ff",x"ff",x"fb",x"f6",x"cd",x"84",x"80",x"80",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"c4",x"a0",x"80",x"80",x"80",x"60",x"60",x"64",x"89",x"b2",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"6e",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"b6",x"ff",x"ff",x"fb",x"d2",x"a9",x"84",x"80",x"a0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e4",x"e4",x"c0",x"c0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"60",x"64",x"89",x"d2",x"f2",x"c9",x"a4",x"a0",x"c0",x"c0",x"e0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"60",x"60",x"64",x"64",x"8d",x"92",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"b6",x"6e",x"6e",x"92",x"db",x"ff",x"ff",x"fb",x"d2",x"89",x"80",x"80",x"a0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"a0",x"80",x"80",x"60",x"40",x"40",x"64",x"8d",x"d6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b2",x"69",x"25",x"49",x"b7",x"ff",x"ff",x"ff",x"f6",x"cd",x"a4",x"80",x"80",x"a0",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"60",x"60",x"64",x"6d",x"b2",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"db",x"b7",x"8e",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"6e",x"d6",x"fb",x"fb",x"f2",x"e9",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c4",x"80",x"60",x"64",x"b2",x"fb",x"ff",x"ff",x"db",x"97",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"6d",x"6d",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"6d",x"db",x"fb",x"b2",x"84",x"60",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a4",x"c9",x"fb",x"ff",x"fb",x"fb",x"f6",x"f6",x"d1",x"cd",x"c9",x"c8",x"c4",x"a4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c4",x"c4",x"e4",x"c9",x"c9",x"e9",x"ed",x"ee",x"f2",x"f2",x"f2",x"f6",x"f6",x"f6",x"f6",x"f6",x"f6",x"d2",x"d2",x"b2",x"d6",x"ff",x"ff",x"b7",x"6e",x"29",x"05",x"05",x"4a",x"b7",x"ff",x"ff",x"fb",x"d6",x"8d",x"84",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"64",x"84",x"89",x"8d",x"b6",x"d7",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"49",x"49",x"8e",x"fb",x"ff",x"ff",x"f7",x"b2",x"a9",x"84",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"60",x"84",x"89",x"8d",x"b2",x"d6",x"db",x"ff",x"ff",x"ff",x"ff",x"df",x"bb",x"6e",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"d7",x"ff",x"ff",x"fb",x"d6",x"ad",x"84",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"60",x"60",x"60",x"64",x"89",x"b2",x"db",x"fb",x"fb",x"d2",x"a5",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"64",x"89",x"8d",x"8d",x"b6",x"db",x"df",x"df",x"ff",x"ff",x"ff",x"ff",x"fb",x"b2",x"69",x"25",x"04",x"04",x"04",x"6e",x"db",x"ff",x"ff",x"ff",x"fb",x"d2",x"ad",x"a9",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"64",x"64",x"89",x"b1",x"b2",x"d6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"49",x"21",x"00",x"00",x"04",x"49",x"96",x"ff",x"ff",x"ff",x"fb",x"f6",x"cd",x"89",x"64",x"60",x"60",x"80",x"80",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"64",x"68",x"89",x"8d",x"b2",x"d6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"4e",x"49",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"49",x"8e",x"d7",x"f7",x"f7",x"f2",x"ed",x"c4",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"60",x"60",x"89",x"d6",x"ff",x"ff",x"ff",x"db",x"92",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"25",x"04",x"00",x"00",x"00",x"24",x"92",x"ff",x"db",x"b2",x"64",x"64",x"84",x"84",x"a4",x"a4",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"a4",x"a4",x"a4",x"c9",x"ed",x"ed",x"f6",x"f6",x"f2",x"ed",x"ed",x"c9",x"c4",x"c4",x"c4",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e5",x"e9",x"e9",x"ed",x"ed",x"f2",x"f2",x"f2",x"f6",x"f6",x"f6",x"f6",x"f6",x"fb",x"fb",x"fb",x"d7",x"b7",x"b2",x"6e",x"6e",x"92",x"d7",x"ff",x"ff",x"ff",x"ff",x"d6",x"b2",x"ad",x"89",x"84",x"84",x"84",x"84",x"84",x"64",x"64",x"64",x"64",x"69",x"8d",x"b2",x"b2",x"d6",x"db",x"df",x"ff",x"ff",x"ff",x"ff",x"fb",x"db",x"b6",x"6e",x"45",x"00",x"00",x"25",x"b2",x"ff",x"ff",x"ff",x"fb",x"d6",x"d2",x"ad",x"a9",x"a4",x"84",x"84",x"84",x"84",x"84",x"80",x"80",x"80",x"60",x"64",x"64",x"64",x"64",x"69",x"8d",x"b2",x"d6",x"db",x"fb",x"ff",x"ff",x"ff",x"ff",x"db",x"b7",x"92",x"6d",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"6e",x"db",x"ff",x"ff",x"fb",x"d6",x"d2",x"ad",x"a9",x"84",x"84",x"84",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"64",x"64",x"64",x"89",x"b2",x"d6",x"fb",x"ff",x"ff",x"ff",x"f7",x"d2",x"a9",x"84",x"84",x"84",x"84",x"84",x"84",x"64",x"68",x"69",x"89",x"8d",x"b2",x"b2",x"b6",x"db",x"df",x"ff",x"ff",x"ff",x"ff",x"db",x"b7",x"b2",x"8e",x"49",x"20",x"00",x"00",x"00",x"00",x"25",x"6e",x"b7",x"ff",x"ff",x"ff",x"ff",x"fb",x"d2",x"ad",x"89",x"84",x"84",x"84",x"84",x"84",x"64",x"64",x"64",x"64",x"64",x"88",x"89",x"89",x"89",x"8d",x"b2",x"d6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b7",x"92",x"6d",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"92",x"db",x"ff",x"ff",x"ff",x"fb",x"b6",x"8d",x"89",x"88",x"84",x"84",x"84",x"84",x"84",x"84",x"64",x"64",x"64",x"64",x"64",x"69",x"89",x"8d",x"b2",x"b6",x"db",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"96",x"6e",x"25",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"49",x"8e",x"b3",x"d7",x"f7",x"f6",x"f2",x"e9",x"e4",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"80",x"60",x"64",x"89",x"b2",x"ff",x"ff",x"ff",x"bb",x"92",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"49",x"d7",x"ff",x"db",x"b6",x"ae",x"ad",x"ad",x"ad",x"b1",x"ad",x"ad",x"b2",x"b1",x"b1",x"ad",x"ad",x"b2",x"b1",x"b1",x"b1",x"ad",x"ad",x"cd",x"cd",x"ed",x"ed",x"f1",x"f1",x"cd",x"e9",x"e5",x"e0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c4",x"c4",x"c4",x"c4",x"e9",x"e9",x"e9",x"ed",x"ed",x"f2",x"f2",x"f6",x"f7",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"d2",x"b2",x"b1",x"ad",x"b2",x"b2",x"b2",x"b6",x"d6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"d7",x"92",x"69",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"92",x"df",x"ff",x"ff",x"ff",x"fb",x"fb",x"f6",x"d2",x"b1",x"8d",x"8d",x"8d",x"69",x"69",x"69",x"69",x"69",x"8d",x"b2",x"b6",x"b6",x"b6",x"d7",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"bb",x"92",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"6e",x"db",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"d6",x"d2",x"b2",x"ad",x"89",x"89",x"89",x"89",x"89",x"89",x"8d",x"ad",x"b2",x"d6",x"db",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"d6",x"b2",x"ad",x"ad",x"ad",x"b2",x"b2",x"b6",x"d6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"ff",x"db",x"92",x"4d",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"4d",x"96",x"df",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"d6",x"d2",x"b2",x"b2",x"b2",x"b1",x"b1",x"b2",x"b2",x"b2",x"b6",x"d6",x"da",x"db",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"92",x"db",x"ff",x"ff",x"ff",x"ff",x"fb",x"db",x"d6",x"d6",x"d2",x"b2",x"b1",x"ad",x"8d",x"8d",x"92",x"b2",x"b2",x"d6",x"d6",x"db",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"69",x"d2",x"fb",x"fb",x"f7",x"f2",x"e9",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"40",x"64",x"ad",x"d6",x"fb",x"ff",x"ff",x"df",x"92",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"4d",x"6d",x"92",x"92",x"92",x"92",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"49",x"24",x"24",x"00",x"00",x"00",x"24",x"b2",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"fb",x"fb",x"fb",x"ff",x"df",x"df",x"df",x"df",x"db",x"fb",x"fb",x"ff",x"ff",x"fb",x"fa",x"f6",x"f6",x"f2",x"ed",x"e9",x"e4",x"c4",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e5",x"e9",x"e9",x"ed",x"f2",x"f2",x"f6",x"f7",x"f7",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"4d",x"29",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"4d",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"bb",x"92",x"4d",x"29",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"49",x"92",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"db",x"d7",x"fb",x"fb",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"bb",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b7",x"92",x"49",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"25",x"6e",x"b7",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b7",x"92",x"4d",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"4d",x"92",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"db",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"db",x"93",x"6e",x"25",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"92",x"b7",x"d7",x"f7",x"f6",x"f2",x"c9",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"89",x"b2",x"fb",x"ff",x"ff",x"ff",x"b7",x"6e",x"25",x"00",x"00",x"00",x"00",x"00",x"04",x"24",x"24",x"49",x"6d",x"71",x"92",x"92",x"92",x"b6",x"b7",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"49",x"24",x"20",x"00",x"00",x"00",x"25",x"b7",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"f6",x"f1",x"ed",x"e9",x"e4",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c4",x"c4",x"e9",x"ed",x"ed",x"ed",x"f1",x"f2",x"f6",x"f6",x"f7",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"92",x"6e",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"92",x"b7",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b7",x"92",x"6d",x"29",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"6e",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b7",x"92",x"6e",x"6e",x"92",x"b7",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"d7",x"b7",x"92",x"8e",x"69",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"49",x"72",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b7",x"92",x"6e",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"29",x"6e",x"92",x"b7",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b7",x"92",x"92",x"6e",x"49",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"25",x"49",x"6e",x"b2",x"d7",x"fb",x"f7",x"f2",x"e9",x"c8",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"60",x"64",x"89",x"b2",x"fb",x"ff",x"ff",x"ff",x"b7",x"6e",x"24",x"00",x"00",x"00",x"00",x"00",x"04",x"24",x"28",x"49",x"49",x"6d",x"92",x"92",x"92",x"b6",x"b7",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"24",x"20",x"00",x"00",x"00",x"29",x"b7",x"db",x"ff",x"ff",x"df",x"df",x"df",x"fb",x"fb",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"f6",x"ee",x"c9",x"c4",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c4",x"c4",x"c4",x"c4",x"c5",x"e9",x"ed",x"ee",x"f2",x"f6",x"fb",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"db",x"b7",x"6e",x"49",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"6d",x"92",x"d7",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"df",x"df",x"db",x"b7",x"92",x"6e",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"49",x"6e",x"92",x"b7",x"db",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"db",x"97",x"6e",x"49",x"25",x"00",x"00",x"25",x"49",x"92",x"b7",x"fb",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"d7",x"b7",x"92",x"6e",x"49",x"25",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"49",x"92",x"b7",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b7",x"b7",x"b7",x"6d",x"49",x"25",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"49",x"6e",x"b3",x"d7",x"db",x"db",x"db",x"df",x"df",x"df",x"ff",x"ff",x"ff",x"db",x"d7",x"b7",x"92",x"8e",x"6e",x"29",x"05",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"45",x"6e",x"92",x"d7",x"fb",x"f7",x"f6",x"f2",x"e9",x"c4",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"40",x"44",x"8d",x"ba",x"ff",x"ff",x"ff",x"ff",x"b7",x"6d",x"24",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"24",x"00",x"00",x"00",x"00",x"05",x"4e",x"6e",x"6e",x"8e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"92",x"b6",x"fb",x"ff",x"ff",x"fb",x"f6",x"f2",x"ee",x"c9",x"c5",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"e0",x"e4",x"e5",x"e9",x"e9",x"ed",x"ed",x"f2",x"f6",x"f6",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"db",x"b7",x"92",x"6e",x"6e",x"49",x"45",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"45",x"49",x"69",x"6e",x"8e",x"92",x"92",x"92",x"92",x"92",x"92",x"72",x"6e",x"6e",x"49",x"49",x"25",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"49",x"49",x"6e",x"72",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6e",x"49",x"49",x"25",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"45",x"49",x"6d",x"6e",x"6e",x"69",x"49",x"49",x"25",x"25",x"25",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"25",x"45",x"49",x"6e",x"6e",x"6e",x"6e",x"6e",x"6d",x"49",x"49",x"49",x"25",x"25",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"25",x"45",x"45",x"49",x"49",x"6d",x"6e",x"6e",x"6e",x"6e",x"49",x"49",x"25",x"25",x"25",x"25",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"6d",x"92",x"b2",x"d7",x"f7",x"f7",x"f2",x"ee",x"c9",x"c4",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"60",x"60",x"89",x"b2",x"db",x"ff",x"ff",x"ff",x"db",x"92",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"49",x"6d",x"8e",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"4d",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"25",x"20",x"20",x"24",x"25",x"05",x"05",x"25",x"25",x"49",x"6e",x"b6",x"fb",x"fb",x"fb",x"f2",x"ed",x"e5",x"e5",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c4",x"c4",x"e9",x"e9",x"ed",x"ed",x"f2",x"f2",x"f6",x"f6",x"f6",x"fb",x"fb",x"fb",x"db",x"d7",x"b6",x"b2",x"8e",x"6d",x"49",x"25",x"25",x"24",x"24",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"25",x"29",x"49",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"25",x"49",x"6d",x"92",x"b6",x"d6",x"fb",x"f7",x"f2",x"ed",x"c9",x"c4",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"64",x"8d",x"d6",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"b6",x"92",x"6d",x"6d",x"4d",x"29",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"49",x"92",x"db",x"ff",x"fb",x"f6",x"ed",x"c5",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e9",x"e9",x"e9",x"cd",x"f1",x"f2",x"f6",x"f6",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"db",x"b7",x"92",x"92",x"6e",x"6d",x"49",x"45",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"49",x"8e",x"b3",x"f7",x"fb",x"fb",x"f6",x"f6",x"f2",x"e9",x"c4",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"40",x"64",x"b2",x"db",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"29",x"04",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"29",x"8e",x"d7",x"fb",x"f7",x"f2",x"cd",x"c9",x"c4",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c4",x"c4",x"e4",x"e9",x"ed",x"cd",x"ed",x"f2",x"f6",x"f6",x"fb",x"fb",x"fb",x"fb",x"db",x"db",x"d7",x"d7",x"b6",x"b2",x"92",x"6e",x"6d",x"49",x"49",x"25",x"05",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"49",x"6e",x"b2",x"d7",x"d7",x"f7",x"f7",x"f2",x"ee",x"ed",x"c9",x"c4",x"c4",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"60",x"89",x"8d",x"b6",x"db",x"ff",x"ff",x"ff",x"bb",x"72",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"6d",x"6d",x"49",x"49",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"29",x"92",x"fb",x"fb",x"f7",x"f2",x"c9",x"a4",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"c0",x"c4",x"c4",x"c4",x"c9",x"c9",x"ed",x"f2",x"f2",x"f6",x"f6",x"f7",x"fb",x"fb",x"fb",x"fb",x"fb",x"db",x"d7",x"b6",x"92",x"92",x"6e",x"49",x"29",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"49",x"49",x"92",x"b6",x"d7",x"fb",x"fb",x"f7",x"f2",x"ee",x"e9",x"c4",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"60",x"60",x"64",x"b2",x"db",x"ff",x"ff",x"df",x"db",x"b7",x"6e",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"6d",x"6d",x"91",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"92",x"db",x"fb",x"fb",x"f2",x"c9",x"c4",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a4",x"a4",x"a4",x"a4",x"a9",x"cd",x"ce",x"f2",x"f6",x"f7",x"fb",x"fb",x"fb",x"fb",x"db",x"db",x"d7",x"d7",x"d7",x"b3",x"b2",x"8e",x"6e",x"49",x"45",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"49",x"6e",x"b2",x"d7",x"fb",x"fb",x"f7",x"f6",x"f2",x"ee",x"cd",x"c9",x"c4",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"64",x"68",x"91",x"d6",x"db",x"ff",x"ff",x"ff",x"db",x"92",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"6d",x"49",x"49",x"25",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"b6",x"fb",x"fb",x"f7",x"f2",x"c9",x"c4",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c4",x"c5",x"c9",x"c9",x"cd",x"cd",x"ce",x"d2",x"d2",x"d6",x"f6",x"f7",x"f7",x"f7",x"f7",x"d7",x"d7",x"b6",x"b2",x"92",x"92",x"72",x"6e",x"6d",x"69",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"49",x"6d",x"92",x"92",x"b6",x"d7",x"d7",x"f7",x"f7",x"f7",x"f2",x"ee",x"e9",x"e9",x"c4",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"60",x"89",x"8d",x"96",x"db",x"ff",x"ff",x"ff",x"ff",x"b6",x"6d",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"91",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"6d",x"49",x"49",x"49",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"25",x"6d",x"b6",x"fb",x"fb",x"f6",x"ed",x"c5",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"84",x"84",x"a5",x"a9",x"a9",x"ce",x"ce",x"ce",x"d2",x"d2",x"d6",x"d6",x"d6",x"d7",x"d7",x"d7",x"d7",x"d6",x"b6",x"b2",x"b2",x"8e",x"6d",x"49",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"49",x"49",x"6d",x"92",x"b7",x"d7",x"fb",x"fb",x"fb",x"f7",x"f6",x"f2",x"ee",x"e9",x"e5",x"e5",x"e0",x"e0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a0",x"80",x"60",x"64",x"69",x"b2",x"db",x"df",x"ff",x"ff",x"ff",x"db",x"b2",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"b2",x"db",x"fb",x"f6",x"ed",x"c4",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"64",x"64",x"84",x"88",x"89",x"8d",x"ad",x"ad",x"ae",x"b2",x"b2",x"d2",x"d6",x"d6",x"b6",x"b2",x"b2",x"b2",x"92",x"92",x"8d",x"69",x"69",x"69",x"49",x"45",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"49",x"6d",x"8e",x"b2",x"b2",x"d6",x"f7",x"fb",x"fb",x"fb",x"f7",x"f7",x"f6",x"f2",x"ed",x"c9",x"c4",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"80",x"60",x"60",x"64",x"8d",x"d2",x"fb",x"fb",x"ff",x"ff",x"ff",x"db",x"b2",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"92",x"fb",x"fb",x"f7",x"cd",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"84",x"84",x"64",x"69",x"89",x"89",x"8d",x"8d",x"8d",x"8d",x"8e",x"b2",x"b2",x"b2",x"b2",x"b2",x"92",x"92",x"92",x"8e",x"6d",x"6d",x"6d",x"4d",x"49",x"49",x"49",x"25",x"25",x"25",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"49",x"49",x"49",x"4d",x"72",x"92",x"92",x"b7",x"db",x"db",x"fb",x"fb",x"f7",x"f7",x"f7",x"f6",x"f2",x"ed",x"ed",x"e9",x"e5",x"c4",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"60",x"64",x"8d",x"b2",x"da",x"ff",x"ff",x"ff",x"ff",x"fb",x"b7",x"6e",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"b7",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"29",x"92",x"db",x"f7",x"f2",x"ed",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"64",x"69",x"69",x"89",x"8d",x"8e",x"8e",x"8e",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6e",x"6e",x"6e",x"69",x"49",x"49",x"25",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"49",x"6d",x"6e",x"92",x"b2",x"b6",x"b6",x"d7",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"f7",x"f6",x"f2",x"ee",x"cd",x"c9",x"c4",x"c4",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"60",x"60",x"44",x"68",x"b1",x"da",x"df",x"df",x"ff",x"ff",x"ff",x"db",x"b2",x"49",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"b7",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"da",x"b6",x"96",x"92",x"6e",x"6d",x"49",x"48",x"44",x"24",x"24",x"00",x"00",x"00",x"00",x"25",x"8e",x"d7",x"fb",x"fb",x"ce",x"c5",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"40",x"64",x"64",x"69",x"69",x"8d",x"8e",x"8e",x"8e",x"8e",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"72",x"72",x"6e",x"6e",x"6d",x"69",x"69",x"49",x"49",x"49",x"29",x"29",x"25",x"25",x"25",x"05",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"05",x"25",x"25",x"29",x"49",x"69",x"6e",x"8e",x"8e",x"92",x"b2",x"b2",x"b6",x"b7",x"db",x"db",x"fb",x"fb",x"fb",x"fb",x"fb",x"f7",x"f7",x"f2",x"f2",x"f2",x"ee",x"ed",x"c9",x"c5",x"c4",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"60",x"40",x"40",x"68",x"8d",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"df",x"b7",x"6e",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"24",x"24",x"28",x"49",x"49",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"d6",x"b6",x"b6",x"92",x"92",x"6e",x"49",x"49",x"44",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"8e",x"d7",x"fb",x"fb",x"f2",x"c5",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"60",x"60",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"40",x"40",x"44",x"64",x"65",x"65",x"69",x"69",x"69",x"69",x"6d",x"6d",x"8d",x"8d",x"8e",x"92",x"92",x"8e",x"8e",x"8e",x"8e",x"8e",x"8e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"69",x"69",x"69",x"49",x"49",x"49",x"49",x"49",x"29",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"04",x"04",x"04",x"00",x"20",x"20",x"20",x"20",x"00",x"00",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"00",x"00",x"04",x"04",x"04",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"6e",x"6e",x"6e",x"72",x"92",x"92",x"92",x"92",x"b2",x"b6",x"d7",x"d7",x"d7",x"f7",x"f7",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"f7",x"f7",x"f2",x"f2",x"ee",x"ee",x"e9",x"e9",x"e5",x"e5",x"c4",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"60",x"64",x"64",x"8d",x"b2",x"da",x"ff",x"ff",x"ff",x"ff",x"ff",x"b7",x"92",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"6d",x"49",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"6d",x"d7",x"fb",x"f7",x"ce",x"c5",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"a4",x"a0",x"80",x"84",x"84",x"84",x"84",x"84",x"80",x"80",x"80",x"84",x"60",x"80",x"80",x"80",x"64",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"64",x"64",x"68",x"69",x"69",x"69",x"69",x"89",x"8d",x"8d",x"8e",x"8e",x"8e",x"8e",x"8e",x"92",x"b2",x"b2",x"b2",x"b2",x"b2",x"92",x"92",x"92",x"92",x"92",x"72",x"72",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6e",x"6e",x"6e",x"8e",x"8e",x"6e",x"6e",x"6d",x"49",x"49",x"49",x"49",x"69",x"6d",x"6d",x"6d",x"4d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"72",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"d7",x"d7",x"d7",x"db",x"db",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"f7",x"f7",x"f7",x"f6",x"f6",x"f2",x"f2",x"f2",x"ee",x"ee",x"ed",x"c9",x"c5",x"c5",x"c5",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"80",x"60",x"60",x"89",x"ad",x"d6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"25",x"6e",x"d7",x"fb",x"f6",x"ed",x"c4",x"c0",x"e0",x"e0",x"e0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"84",x"84",x"84",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"c4",x"c4",x"a4",x"c4",x"c4",x"c4",x"c4",x"c4",x"c8",x"c8",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c8",x"c8",x"c8",x"a8",x"c8",x"c8",x"c8",x"e8",x"e8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"e8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"a8",x"a8",x"c4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"44",x"44",x"64",x"64",x"64",x"68",x"69",x"69",x"6d",x"6d",x"6d",x"8e",x"92",x"92",x"92",x"b2",x"b2",x"b2",x"d2",x"d2",x"d6",x"d6",x"d6",x"d6",x"d7",x"d7",x"d7",x"d7",x"d7",x"d7",x"d7",x"d7",x"db",x"fb",x"fb",x"fb",x"db",x"d7",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"f7",x"f7",x"f7",x"f7",x"f7",x"f7",x"f7",x"f7",x"f7",x"f2",x"f2",x"f2",x"f2",x"ee",x"ee",x"ed",x"ed",x"e9",x"e9",x"c9",x"c9",x"c5",x"e4",x"e4",x"e0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"60",x"64",x"69",x"8d",x"b2",x"d6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"b7",x"92",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"72",x"6d",x"6d",x"6d",x"49",x"24",x"20",x"00",x"00",x"00",x"00",x"04",x"6e",x"b7",x"fb",x"f6",x"ed",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"84",x"a4",x"a4",x"a4",x"a4",x"a4",x"c8",x"c8",x"c8",x"e8",x"e8",x"e8",x"e8",x"c8",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c8",x"c8",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"c4",x"a4",x"a4",x"a4",x"a4",x"84",x"84",x"84",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"44",x"44",x"45",x"65",x"69",x"69",x"89",x"89",x"89",x"89",x"a9",x"ad",x"ad",x"ad",x"ad",x"ad",x"ae",x"ae",x"ce",x"d2",x"d2",x"d2",x"d2",x"f2",x"f6",x"f6",x"f6",x"f6",x"f6",x"f6",x"f6",x"f6",x"f7",x"f7",x"f7",x"f7",x"f7",x"f7",x"f7",x"f7",x"f7",x"f7",x"f7",x"f7",x"f7",x"f7",x"f7",x"f7",x"f7",x"f6",x"f6",x"f7",x"f2",x"f2",x"f2",x"f2",x"f2",x"ee",x"ee",x"ee",x"ee",x"ed",x"ed",x"ed",x"e9",x"e9",x"e5",x"e5",x"e5",x"e5",x"e5",x"e4",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"64",x"68",x"8d",x"b6",x"bb",x"df",x"ff",x"ff",x"ff",x"ff",x"db",x"b7",x"92",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"6d",x"6d",x"6d",x"49",x"45",x"24",x"00",x"00",x"00",x"00",x"00",x"4e",x"d7",x"fb",x"f7",x"ce",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"60",x"60",x"80",x"80",x"80",x"80",x"84",x"a4",x"a4",x"a4",x"c8",x"c8",x"c8",x"c8",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"c8",x"c8",x"c8",x"c8",x"c8",x"c8",x"e8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"e8",x"c8",x"c8",x"c4",x"a4",x"a4",x"a0",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"84",x"84",x"84",x"a4",x"a4",x"a4",x"a4",x"c9",x"c9",x"c9",x"c9",x"c9",x"c9",x"e9",x"e9",x"e9",x"e9",x"c9",x"c9",x"c9",x"c9",x"c9",x"c9",x"c9",x"c5",x"c5",x"c5",x"c5",x"c5",x"c5",x"c5",x"c5",x"c4",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"60",x"60",x"64",x"8d",x"b2",x"d6",x"db",x"ff",x"ff",x"ff",x"ff",x"df",x"db",x"b7",x"6e",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"4d",x"49",x"44",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"b7",x"fb",x"fb",x"cd",x"c5",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"84",x"84",x"a4",x"a4",x"c4",x"c4",x"c4",x"c8",x"c8",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"c4",x"c4",x"c8",x"c4",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"c8",x"c8",x"cd",x"d1",x"d1",x"d1",x"cd",x"cd",x"ed",x"e8",x"e8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c8",x"c8",x"cd",x"cd",x"cd",x"cd",x"c8",x"c8",x"c8",x"e8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"c4",x"c4",x"c4",x"a4",x"a4",x"a4",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"60",x"60",x"60",x"64",x"89",x"b2",x"d6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"bb",x"92",x"4d",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"92",x"92",x"92",x"4d",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"b2",x"fb",x"fb",x"f2",x"a4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"a4",x"a4",x"a4",x"c8",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c8",x"c8",x"c8",x"cc",x"cc",x"c8",x"c8",x"e4",x"e4",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"c8",x"c4",x"c8",x"cc",x"d1",x"f6",x"f6",x"fa",x"fa",x"fa",x"f6",x"f2",x"f1",x"ed",x"e8",x"e4",x"e4",x"e4",x"e4",x"c8",x"c8",x"cc",x"d1",x"d1",x"d6",x"d6",x"f6",x"f6",x"f1",x"f1",x"cc",x"e8",x"e4",x"e4",x"e8",x"e8",x"e8",x"c8",x"c8",x"c8",x"c8",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c8",x"c4",x"c4",x"c4",x"a4",x"a0",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"60",x"64",x"64",x"68",x"8d",x"b2",x"d6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b7",x"92",x"6d",x"29",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"48",x"48",x"48",x"48",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"4d",x"49",x"24",x"20",x"00",x"00",x"00",x"00",x"25",x"b2",x"fb",x"f7",x"ed",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"64",x"64",x"64",x"68",x"68",x"68",x"68",x"68",x"69",x"69",x"89",x"89",x"69",x"64",x"64",x"64",x"64",x"64",x"64",x"64",x"64",x"64",x"64",x"64",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"a0",x"a4",x"a4",x"c4",x"c8",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"c8",x"c8",x"ed",x"f1",x"f6",x"f6",x"f1",x"ed",x"e8",x"e4",x"e4",x"e4",x"e8",x"e4",x"e4",x"e4",x"c4",x"c8",x"cd",x"f6",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fa",x"f6",x"ed",x"e4",x"e4",x"e4",x"c4",x"c8",x"d1",x"d6",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fa",x"f6",x"ed",x"e8",x"e4",x"e4",x"e4",x"c8",x"cc",x"d1",x"d1",x"f1",x"ed",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"c4",x"c4",x"c8",x"a8",x"c8",x"c8",x"c8",x"c8",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"c4",x"c4",x"c4",x"a4",x"a4",x"84",x"80",x"60",x"60",x"60",x"60",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"80",x"60",x"60",x"60",x"64",x"8d",x"b1",x"b6",x"da",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"6e",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"48",x"49",x"49",x"69",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"25",x"6e",x"fb",x"fb",x"f2",x"c4",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"84",x"84",x"84",x"89",x"a9",x"a9",x"ad",x"ad",x"ad",x"ad",x"b2",x"b6",x"b6",x"b6",x"b6",x"d6",x"d6",x"d6",x"d6",x"d6",x"d6",x"d6",x"d6",x"d6",x"d6",x"d6",x"d6",x"d6",x"d6",x"b6",x"b2",x"b2",x"b2",x"b2",x"b2",x"b1",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"a9",x"a9",x"a9",x"a9",x"a9",x"a9",x"a4",x"84",x"84",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"a4",x"a4",x"c4",x"c4",x"e4",x"e4",x"e4",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"c8",x"c8",x"a8",x"c8",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"c8",x"f1",x"f6",x"fb",x"ff",x"ff",x"fa",x"f2",x"ed",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"c4",x"cd",x"f6",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"f6",x"ed",x"e4",x"e4",x"e4",x"c4",x"cd",x"d6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fa",x"f1",x"e8",x"e4",x"e4",x"c4",x"e8",x"f1",x"fa",x"fa",x"fa",x"f2",x"e9",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"c4",x"c8",x"c8",x"cd",x"cd",x"d1",x"d1",x"cd",x"cc",x"cc",x"c8",x"c8",x"c8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"c8",x"c4",x"c4",x"c4",x"a4",x"a4",x"a4",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"64",x"84",x"89",x"ad",x"b2",x"d6",x"db",x"df",x"ff",x"ff",x"ff",x"ff",x"df",x"bb",x"96",x"72",x"49",x"45",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"6d",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"4d",x"d7",x"fb",x"f6",x"c9",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"64",x"64",x"64",x"69",x"8d",x"8d",x"b2",x"d6",x"d6",x"d6",x"db",x"fb",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"fb",x"fb",x"fb",x"db",x"d6",x"d6",x"d6",x"d6",x"d6",x"d6",x"b2",x"ad",x"ad",x"8d",x"89",x"89",x"64",x"64",x"64",x"84",x"84",x"84",x"84",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a4",x"c4",x"c4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"c8",x"c8",x"cc",x"ad",x"cc",x"c8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"ed",x"f6",x"ff",x"ff",x"ff",x"ff",x"ff",x"f6",x"ed",x"c4",x"c4",x"e4",x"e4",x"e4",x"e0",x"c0",x"c4",x"f2",x"fb",x"ff",x"ff",x"ff",x"fb",x"f6",x"f6",x"f6",x"fb",x"ff",x"fa",x"f5",x"ed",x"c4",x"e4",x"e4",x"e8",x"f2",x"fb",x"ff",x"ff",x"ff",x"fb",x"fa",x"fa",x"ff",x"ff",x"ff",x"fb",x"f2",x"e9",x"e4",x"e4",x"e4",x"e9",x"f6",x"ff",x"ff",x"ff",x"f6",x"ed",x"c4",x"e4",x"e4",x"e4",x"c4",x"c4",x"c8",x"c9",x"cd",x"f2",x"f6",x"f6",x"fa",x"fa",x"f6",x"f6",x"f5",x"d1",x"cd",x"c8",x"c4",x"c4",x"e4",x"e4",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"a4",x"a4",x"a4",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"64",x"64",x"64",x"8d",x"b2",x"d6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"92",x"6e",x"29",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"44",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6e",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"29",x"b7",x"ff",x"f6",x"cd",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a0",x"80",x"80",x"60",x"64",x"64",x"89",x"91",x"b2",x"b6",x"bb",x"db",x"db",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"fb",x"fb",x"d6",x"d6",x"d6",x"d2",x"b1",x"ad",x"ad",x"ad",x"a9",x"a9",x"88",x"84",x"84",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"a4",x"a4",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"c4",x"c4",x"c4",x"c8",x"c8",x"cc",x"cd",x"ed",x"ed",x"ed",x"ed",x"c4",x"c4",x"c4",x"c4",x"c8",x"f1",x"fa",x"fa",x"fa",x"f1",x"c8",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c8",x"f2",x"fb",x"ff",x"ff",x"df",x"df",x"ff",x"fb",x"f2",x"c8",x"c4",x"e4",x"e4",x"e0",x"e0",x"c0",x"c4",x"f6",x"ff",x"ff",x"ff",x"fb",x"d2",x"ed",x"e9",x"e9",x"f1",x"f6",x"f5",x"cd",x"c8",x"c4",x"c4",x"e8",x"ed",x"f6",x"ff",x"ff",x"ff",x"fa",x"d2",x"cd",x"cd",x"d2",x"f6",x"fb",x"fb",x"f2",x"c4",x"e4",x"e4",x"e0",x"e9",x"f6",x"ff",x"ff",x"ff",x"f6",x"ed",x"e4",x"e4",x"e4",x"c4",x"c4",x"c8",x"cd",x"f2",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f2",x"ed",x"c8",x"c4",x"e4",x"e4",x"e4",x"e4",x"c8",x"c8",x"c4",x"c4",x"c4",x"c4",x"c4",x"c4",x"c4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c8",x"c4",x"c4",x"a4",x"a0",x"80",x"80",x"80",x"80",x"a0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"64",x"89",x"8d",x"b6",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"db",x"92",x"6e",x"25",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6e",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"20",x"00",x"00",x"00",x"00",x"92",x"fb",x"fb",x"ee",x"c5",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"60",x"40",x"60",x"84",x"89",x"ad",x"b2",x"b2",x"d6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b6",x"b6",x"b6",x"b6",x"b6",x"96",x"96",x"b6",x"b7",x"b7",x"b7",x"b7",x"b7",x"bb",x"db",x"db",x"db",x"db",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"db",x"db",x"db",x"d6",x"d6",x"d6",x"d2",x"b2",x"ad",x"ad",x"ad",x"a9",x"a9",x"a9",x"a5",x"84",x"84",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"c0",x"a0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"60",x"80",x"c4",x"c4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e4",x"e8",x"e4",x"e4",x"e4",x"c4",x"a8",x"cd",x"d1",x"d2",x"f6",x"fa",x"fa",x"fa",x"fa",x"f6",x"f1",x"c9",x"a4",x"c4",x"cd",x"f6",x"ff",x"ff",x"ff",x"f6",x"e9",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e4",x"c9",x"f6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"f6",x"c9",x"c0",x"e4",x"e4",x"e0",x"e0",x"c4",x"c9",x"f6",x"ff",x"ff",x"ff",x"f6",x"cd",x"c4",x"c0",x"c4",x"e8",x"e8",x"e8",x"c8",x"c4",x"c4",x"c4",x"c8",x"f1",x"fb",x"ff",x"ff",x"fb",x"f6",x"c9",x"a4",x"c4",x"c8",x"e9",x"ed",x"ed",x"e9",x"e4",x"e4",x"e4",x"e0",x"e9",x"f6",x"ff",x"ff",x"ff",x"fa",x"ed",x"e4",x"e4",x"e4",x"e4",x"c4",x"cd",x"f6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"f1",x"c8",x"c4",x"e4",x"e4",x"c4",x"a8",x"cd",x"d1",x"d1",x"f2",x"f1",x"cd",x"cd",x"c8",x"c8",x"c4",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"c4",x"80",x"60",x"60",x"80",x"80",x"a0",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"60",x"64",x"84",x"89",x"8d",x"8d",x"b2",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"6d",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"49",x"d7",x"fb",x"f2",x"e9",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"60",x"60",x"44",x"44",x"6d",x"92",x"d6",x"db",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"db",x"db",x"db",x"b7",x"b7",x"b6",x"92",x"92",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"92",x"92",x"92",x"92",x"b6",x"b7",x"b7",x"b7",x"db",x"db",x"db",x"db",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"db",x"db",x"d7",x"d6",x"d6",x"b2",x"b2",x"8d",x"89",x"89",x"64",x"64",x"64",x"64",x"64",x"84",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"80",x"80",x"60",x"60",x"80",x"e4",x"e4",x"e4",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"c8",x"cd",x"d6",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d1",x"c4",x"c4",x"ed",x"fa",x"ff",x"ff",x"ff",x"f2",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e4",x"e4",x"e4",x"e4",x"e0",x"c4",x"cd",x"fb",x"ff",x"ff",x"fb",x"ff",x"ff",x"ff",x"ff",x"fb",x"cd",x"c4",x"c4",x"e4",x"e4",x"e0",x"c4",x"c9",x"f6",x"ff",x"ff",x"ff",x"f6",x"cd",x"a4",x"a0",x"a0",x"c4",x"e4",x"e4",x"c4",x"c4",x"e4",x"c4",x"c4",x"f1",x"fb",x"ff",x"ff",x"ff",x"f6",x"c9",x"c4",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"c0",x"c9",x"f6",x"ff",x"ff",x"ff",x"fa",x"ed",x"e4",x"e4",x"e4",x"c4",x"e9",x"f2",x"fb",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"f6",x"c8",x"c4",x"c0",x"c4",x"c8",x"ad",x"d6",x"fa",x"fb",x"ff",x"ff",x"f6",x"f6",x"f1",x"cd",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"80",x"60",x"60",x"80",x"80",x"80",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"64",x"69",x"8d",x"b2",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"db",x"db",x"b6",x"92",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"49",x"b7",x"fb",x"f2",x"c9",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"60",x"64",x"89",x"b1",x"d6",x"db",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b7",x"92",x"6e",x"6d",x"49",x"25",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b7",x"db",x"db",x"db",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"fa",x"f6",x"d6",x"b2",x"b1",x"8d",x"8d",x"89",x"68",x"64",x"64",x"64",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"60",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"c4",x"c4",x"cc",x"d1",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f1",x"c4",x"c4",x"ed",x"f6",x"ff",x"ff",x"ff",x"f2",x"e8",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"c8",x"d6",x"ff",x"ff",x"ff",x"d6",x"d6",x"fb",x"ff",x"ff",x"ff",x"f6",x"c9",x"c0",x"e0",x"e4",x"e4",x"e4",x"cd",x"fa",x"ff",x"ff",x"ff",x"ff",x"fa",x"d1",x"c9",x"c8",x"c4",x"c0",x"c0",x"e4",x"e4",x"e4",x"e0",x"e4",x"ed",x"f6",x"fb",x"ff",x"ff",x"ff",x"d2",x"c9",x"c4",x"c0",x"c0",x"c0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"c9",x"f6",x"ff",x"ff",x"ff",x"fa",x"cd",x"c4",x"e4",x"c4",x"c4",x"ed",x"f6",x"ff",x"ff",x"ff",x"fb",x"f6",x"f2",x"ee",x"cd",x"cd",x"d6",x"f6",x"fb",x"ff",x"fb",x"f6",x"e9",x"c4",x"c4",x"e8",x"f1",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fa",x"f1",x"e9",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"80",x"60",x"60",x"80",x"80",x"80",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"a0",x"80",x"60",x"60",x"60",x"60",x"64",x"84",x"89",x"ad",x"b2",x"b2",x"d6",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b7",x"92",x"6d",x"49",x"45",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"72",x"fb",x"f7",x"ee",x"c4",x"c0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"65",x"89",x"91",x"b6",x"da",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b7",x"92",x"6e",x"4d",x"49",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"25",x"25",x"49",x"49",x"49",x"69",x"6d",x"6e",x"72",x"92",x"92",x"b6",x"b7",x"b7",x"db",x"db",x"db",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"db",x"db",x"da",x"d6",x"b6",x"b2",x"b2",x"8d",x"8d",x"8d",x"89",x"88",x"84",x"84",x"84",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"20",x"20",x"60",x"c4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e4",x"e4",x"c4",x"c4",x"c8",x"d5",x"fa",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"fb",x"ff",x"ff",x"ff",x"f6",x"ed",x"e4",x"c4",x"ed",x"fa",x"ff",x"ff",x"ff",x"f2",x"e8",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e0",x"e4",x"e4",x"e4",x"e0",x"e4",x"c4",x"cd",x"fa",x"ff",x"ff",x"ff",x"d1",x"cd",x"f6",x"ff",x"ff",x"ff",x"fa",x"d1",x"e4",x"e0",x"e4",x"e0",x"c4",x"c8",x"f2",x"fb",x"ff",x"ff",x"ff",x"ff",x"fa",x"d6",x"d1",x"cd",x"c4",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"ed",x"f6",x"fb",x"ff",x"ff",x"ff",x"fb",x"f6",x"f2",x"c9",x"c4",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"ed",x"f6",x"ff",x"ff",x"ff",x"fa",x"cd",x"c0",x"c4",x"c4",x"c8",x"f6",x"fb",x"ff",x"ff",x"ff",x"f6",x"cd",x"c9",x"c4",x"c4",x"c4",x"c9",x"ed",x"f2",x"f6",x"f6",x"f1",x"e4",x"c0",x"c4",x"ed",x"f6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fa",x"f1",x"c4",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"80",x"60",x"60",x"80",x"80",x"80",x"a0",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"64",x"64",x"68",x"89",x"8d",x"8d",x"b2",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b7",x"92",x"6e",x"49",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"49",x"b6",x"fb",x"f2",x"c9",x"c0",x"c0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"60",x"64",x"89",x"b2",x"d7",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b7",x"92",x"6e",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"49",x"49",x"6d",x"6e",x"6e",x"92",x"92",x"b2",x"b7",x"bb",x"bb",x"bb",x"bb",x"df",x"df",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"fb",x"d7",x"d6",x"b2",x"92",x"92",x"8d",x"89",x"69",x"64",x"44",x"40",x"20",x"20",x"20",x"20",x"60",x"c4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"c4",x"a4",x"c8",x"d1",x"da",x"ff",x"ff",x"ff",x"fb",x"f6",x"f2",x"f2",x"f2",x"f6",x"fa",x"f6",x"f1",x"e8",x"e4",x"c4",x"ed",x"fa",x"ff",x"ff",x"ff",x"f2",x"e8",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"c0",x"c4",x"d1",x"ff",x"ff",x"ff",x"fb",x"c9",x"c9",x"f2",x"fb",x"ff",x"ff",x"ff",x"d6",x"e4",x"e4",x"e4",x"e0",x"c0",x"c4",x"ed",x"f2",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"da",x"d2",x"cd",x"c9",x"c4",x"c0",x"e0",x"e0",x"e0",x"e8",x"ed",x"f6",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"d1",x"cd",x"c8",x"c4",x"c0",x"e0",x"e0",x"e0",x"e9",x"f6",x"ff",x"ff",x"ff",x"fa",x"cd",x"c0",x"c0",x"c4",x"cd",x"fa",x"ff",x"ff",x"ff",x"fb",x"f1",x"c8",x"c4",x"c0",x"c0",x"c0",x"c4",x"c4",x"e9",x"ed",x"ed",x"e9",x"e4",x"c0",x"c4",x"ed",x"f6",x"ff",x"ff",x"ff",x"fb",x"f6",x"f6",x"fb",x"ff",x"ff",x"ff",x"ff",x"f2",x"c0",x"c0",x"e0",x"e4",x"e4",x"e4",x"e4",x"c4",x"80",x"60",x"60",x"80",x"80",x"80",x"a0",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"69",x"8d",x"92",x"b6",x"d6",x"da",x"db",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b7",x"92",x"8e",x"69",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"b7",x"fb",x"f7",x"c9",x"c4",x"c0",x"e4",x"c0",x"80",x"60",x"60",x"85",x"8d",x"b1",x"d6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b7",x"92",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"04",x"00",x"00",x"00",x"00",x"04",x"04",x"04",x"04",x"04",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"04",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"25",x"25",x"49",x"4d",x"6e",x"92",x"96",x"b7",x"b7",x"db",x"db",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"db",x"d7",x"b6",x"92",x"8d",x"69",x"49",x"49",x"44",x"64",x"c4",x"e4",x"e0",x"e4",x"e0",x"e0",x"e0",x"c4",x"a8",x"f1",x"fa",x"ff",x"ff",x"ff",x"f6",x"ed",x"c9",x"c4",x"c4",x"c4",x"c4",x"c5",x"c4",x"e8",x"e4",x"e0",x"c4",x"ed",x"fa",x"ff",x"ff",x"ff",x"f2",x"e9",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"c0",x"c9",x"f6",x"ff",x"ff",x"fb",x"f2",x"c4",x"c4",x"ed",x"f6",x"ff",x"ff",x"ff",x"f6",x"e4",x"e0",x"e4",x"e0",x"e0",x"e0",x"e4",x"e9",x"f2",x"f7",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"cd",x"c9",x"e4",x"e0",x"e0",x"c4",x"c4",x"cd",x"f6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fa",x"d1",x"c9",x"c4",x"c0",x"e0",x"e0",x"e9",x"f6",x"ff",x"ff",x"ff",x"fa",x"ed",x"c0",x"e0",x"e4",x"ed",x"fb",x"ff",x"ff",x"ff",x"f6",x"c9",x"c4",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"c0",x"c0",x"c0",x"ed",x"fb",x"ff",x"ff",x"ff",x"f6",x"a9",x"a4",x"a9",x"cd",x"f6",x"fa",x"f6",x"f1",x"c0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"c0",x"80",x"60",x"40",x"60",x"80",x"80",x"a0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"84",x"84",x"89",x"a9",x"ad",x"b2",x"b2",x"d6",x"d6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"db",x"b7",x"92",x"6e",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"49",x"db",x"fb",x"f2",x"c4",x"a0",x"c0",x"a0",x"80",x"60",x"64",x"69",x"b2",x"d6",x"db",x"ff",x"ff",x"ff",x"ff",x"db",x"d7",x"b3",x"6e",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"25",x"49",x"49",x"49",x"6e",x"6e",x"92",x"92",x"b6",x"b7",x"b7",x"db",x"db",x"db",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"db",x"b6",x"92",x"92",x"6e",x"69",x"84",x"c4",x"e4",x"e0",x"e4",x"e0",x"e0",x"c0",x"c4",x"cd",x"f6",x"ff",x"ff",x"ff",x"f6",x"ed",x"e4",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"c4",x"ed",x"fa",x"ff",x"ff",x"ff",x"f2",x"e8",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"c4",x"d1",x"fa",x"ff",x"ff",x"f7",x"cd",x"a0",x"a0",x"c8",x"f2",x"fb",x"ff",x"ff",x"fb",x"e9",x"c4",x"c0",x"e4",x"e0",x"e0",x"e0",x"e4",x"e9",x"ed",x"f2",x"f6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"fa",x"d1",x"e8",x"e0",x"e0",x"c4",x"c4",x"c4",x"e9",x"f1",x"f6",x"fa",x"fb",x"ff",x"ff",x"ff",x"ff",x"fb",x"f2",x"c8",x"c4",x"e0",x"e0",x"e9",x"f6",x"ff",x"ff",x"ff",x"fa",x"ed",x"c0",x"e0",x"e4",x"ee",x"fb",x"ff",x"ff",x"ff",x"f6",x"c8",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"ed",x"fb",x"ff",x"ff",x"ff",x"f6",x"c9",x"a0",x"a0",x"c4",x"c9",x"ed",x"ed",x"e8",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"c0",x"80",x"40",x"40",x"60",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"84",x"84",x"84",x"89",x"89",x"89",x"8d",x"b2",x"b2",x"d6",x"d6",x"db",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"db",x"d7",x"b2",x"92",x"6e",x"49",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"24",x"24",x"00",x"00",x"00",x"45",x"92",x"fb",x"f7",x"ed",x"a0",x"a0",x"a0",x"60",x"60",x"69",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"df",x"b7",x"92",x"6a",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"28",x"29",x"28",x"24",x"24",x"24",x"24",x"28",x"48",x"48",x"48",x"48",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"49",x"49",x"49",x"44",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"24",x"25",x"29",x"49",x"49",x"4d",x"6e",x"72",x"92",x"96",x"b6",x"bb",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"bb",x"b6",x"96",x"96",x"6d",x"89",x"c9",x"e4",x"e0",x"e0",x"e0",x"e0",x"c0",x"c4",x"cd",x"fb",x"ff",x"ff",x"fa",x"f1",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"ed",x"fb",x"ff",x"ff",x"ff",x"f2",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"c0",x"c4",x"f6",x"ff",x"ff",x"ff",x"f6",x"a9",x"84",x"80",x"a8",x"d2",x"fb",x"fb",x"ff",x"ff",x"f2",x"c5",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c4",x"c4",x"c8",x"ed",x"f6",x"fb",x"ff",x"ff",x"ff",x"ff",x"fa",x"c8",x"c0",x"e0",x"e4",x"e4",x"e0",x"c0",x"c4",x"e9",x"ed",x"f6",x"fb",x"ff",x"ff",x"ff",x"ff",x"fb",x"ed",x"c4",x"e0",x"e0",x"c8",x"d6",x"ff",x"ff",x"ff",x"fa",x"ed",x"c0",x"c0",x"e4",x"f2",x"fb",x"ff",x"ff",x"ff",x"f2",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"ed",x"f6",x"ff",x"ff",x"ff",x"fb",x"ed",x"c4",x"c0",x"c0",x"c0",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"c4",x"80",x"40",x"40",x"60",x"80",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"64",x"89",x"8d",x"b2",x"d6",x"d6",x"d6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"d7",x"b7",x"92",x"8e",x"69",x"45",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"49",x"49",x"24",x"00",x"00",x"00",x"20",x"8e",x"db",x"fb",x"d2",x"a5",x"80",x"60",x"80",x"84",x"8d",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"bb",x"92",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"4d",x"6d",x"6d",x"6d",x"4d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"25",x"25",x"25",x"45",x"49",x"49",x"4d",x"6d",x"6e",x"6e",x"6e",x"6e",x"69",x"64",x"c5",x"e4",x"e0",x"e0",x"e0",x"e0",x"c0",x"c9",x"f6",x"ff",x"ff",x"ff",x"d6",x"c9",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"ed",x"fb",x"ff",x"ff",x"ff",x"f2",x"e4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"c0",x"c4",x"cd",x"fa",x"ff",x"ff",x"ff",x"f7",x"d2",x"ad",x"ad",x"d1",x"d6",x"fb",x"ff",x"ff",x"ff",x"f7",x"cd",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e0",x"c0",x"c0",x"e0",x"e5",x"ee",x"fb",x"ff",x"df",x"ff",x"fa",x"c9",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c4",x"cd",x"f6",x"ff",x"ff",x"ff",x"fb",x"f2",x"e8",x"e0",x"e0",x"c8",x"d6",x"ff",x"ff",x"ff",x"fa",x"cd",x"c0",x"c0",x"c4",x"f2",x"fb",x"ff",x"ff",x"ff",x"f2",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c4",x"ed",x"fb",x"ff",x"ff",x"ff",x"fa",x"f1",x"c4",x"c0",x"c0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e4",x"c0",x"60",x"40",x"40",x"40",x"60",x"60",x"80",x"80",x"80",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"64",x"64",x"84",x"89",x"89",x"8d",x"ad",x"b2",x"b2",x"b2",x"d6",x"d6",x"d6",x"db",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b7",x"b7",x"92",x"6e",x"49",x"25",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"92",x"6d",x"6d",x"49",x"24",x"00",x"00",x"00",x"00",x"45",x"b7",x"fb",x"d2",x"a9",x"60",x"60",x"64",x"88",x"b2",x"db",x"df",x"ff",x"ff",x"ff",x"db",x"b6",x"6e",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"44",x"44",x"44",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"48",x"48",x"28",x"28",x"28",x"24",x"24",x"24",x"24",x"24",x"24",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"24",x"24",x"25",x"25",x"24",x"60",x"a4",x"e4",x"e0",x"e0",x"e0",x"e0",x"c4",x"cd",x"fb",x"ff",x"ff",x"ff",x"d2",x"c8",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c9",x"fb",x"ff",x"ff",x"ff",x"f2",x"e8",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c8",x"f2",x"fb",x"ff",x"ff",x"ff",x"fb",x"d7",x"d6",x"d6",x"fa",x"fb",x"ff",x"ff",x"ff",x"ff",x"fb",x"f2",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e4",x"c0",x"c0",x"c0",x"c0",x"c0",x"c9",x"f6",x"ff",x"ff",x"ff",x"fa",x"c9",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a4",x"d2",x"fb",x"ff",x"ff",x"fb",x"f6",x"e9",x"e0",x"e0",x"c9",x"d6",x"ff",x"ff",x"ff",x"fa",x"cd",x"c0",x"c0",x"c4",x"cd",x"fb",x"ff",x"ff",x"ff",x"f2",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e0",x"e0",x"e0",x"e0",x"e4",x"e0",x"e0",x"e0",x"c0",x"c9",x"f2",x"fa",x"ff",x"ff",x"ff",x"fa",x"f2",x"c9",x"c4",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"60",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"84",x"84",x"84",x"89",x"89",x"89",x"8d",x"8d",x"b1",x"b2",x"b6",x"b6",x"d6",x"db",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"df",x"db",x"bb",x"b7",x"b7",x"92",x"92",x"6e",x"69",x"49",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"48",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"6d",x"6d",x"49",x"24",x"00",x"00",x"00",x"00",x"6e",x"db",x"fb",x"8d",x"64",x"40",x"89",x"ad",x"b2",x"db",x"ff",x"ff",x"ff",x"db",x"b6",x"6d",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"69",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"8e",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"48",x"29",x"29",x"29",x"24",x"24",x"24",x"24",x"04",x"04",x"04",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"a4",x"e4",x"e0",x"e0",x"e0",x"e0",x"c4",x"f2",x"fb",x"ff",x"ff",x"fb",x"cd",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c9",x"fb",x"ff",x"ff",x"ff",x"f2",x"e9",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"a4",x"cd",x"f6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"cd",x"c0",x"c0",x"c0",x"c4",x"c4",x"a4",x"a4",x"a4",x"c0",x"c0",x"a0",x"a9",x"f6",x"ff",x"ff",x"ff",x"fa",x"e9",x"e0",x"e0",x"c0",x"c0",x"c4",x"c4",x"c4",x"c4",x"a0",x"a0",x"80",x"ad",x"f7",x"ff",x"ff",x"ff",x"fa",x"e9",x"c0",x"e0",x"c9",x"d6",x"ff",x"ff",x"ff",x"fa",x"cd",x"c0",x"e0",x"e4",x"c9",x"f6",x"ff",x"ff",x"ff",x"f6",x"c9",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c4",x"e9",x"f2",x"f6",x"fb",x"ff",x"ff",x"fb",x"f6",x"f1",x"c9",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"40",x"20",x"00",x"20",x"00",x"00",x"20",x"40",x"44",x"64",x"64",x"69",x"69",x"8d",x"8d",x"8d",x"b2",x"b6",x"b6",x"d6",x"d6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"df",x"db",x"b7",x"96",x"92",x"72",x"6e",x"49",x"49",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"4d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"24",x"00",x"00",x"00",x"20",x"b3",x"fb",x"d6",x"44",x"44",x"8d",x"b6",x"db",x"df",x"ff",x"ff",x"df",x"b7",x"6e",x"29",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"4d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6e",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"69",x"49",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"44",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"a4",x"e4",x"e0",x"e4",x"e0",x"c0",x"c8",x"f2",x"ff",x"ff",x"ff",x"f7",x"ed",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"cd",x"fb",x"ff",x"ff",x"ff",x"f2",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a4",x"d1",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"ed",x"a0",x"c0",x"c4",x"ed",x"f2",x"f2",x"f1",x"ed",x"c9",x"c8",x"cd",x"d2",x"fb",x"ff",x"ff",x"ff",x"f7",x"e9",x"c0",x"c0",x"e8",x"ed",x"f2",x"f6",x"f1",x"c8",x"a4",x"a4",x"85",x"b2",x"fb",x"ff",x"ff",x"ff",x"fa",x"c9",x"c0",x"e0",x"c9",x"d6",x"ff",x"ff",x"ff",x"fb",x"ed",x"c0",x"e0",x"e0",x"c4",x"f6",x"ff",x"ff",x"ff",x"fb",x"f2",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e9",x"f2",x"f6",x"fb",x"ff",x"ff",x"ff",x"fb",x"f6",x"ed",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"a4",x"64",x"24",x"24",x"44",x"49",x"4d",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"bb",x"db",x"db",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"db",x"db",x"b7",x"b6",x"92",x"6e",x"69",x"49",x"49",x"25",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"48",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"71",x"92",x"92",x"92",x"92",x"92",x"b2",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"49",x"24",x"00",x"00",x"00",x"00",x"49",x"db",x"db",x"b2",x"69",x"8d",x"d6",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"49",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"4d",x"6d",x"6d",x"6d",x"6d",x"72",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"49",x"49",x"49",x"48",x"44",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"a4",x"e0",x"e0",x"e4",x"e0",x"c0",x"c4",x"f2",x"ff",x"ff",x"ff",x"fb",x"cd",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"e0",x"e0",x"c0",x"ed",x"fb",x"ff",x"ff",x"ff",x"f2",x"c4",x"a0",x"c0",x"e0",x"e4",x"e4",x"e0",x"e0",x"c0",x"c0",x"c8",x"d6",x"ff",x"ff",x"ff",x"ff",x"d6",x"f6",x"f7",x"f6",x"f6",x"f6",x"f6",x"f6",x"fb",x"ff",x"ff",x"ff",x"fb",x"f2",x"a4",x"a0",x"c9",x"f6",x"fb",x"fb",x"fb",x"f6",x"f2",x"f2",x"f6",x"fb",x"ff",x"ff",x"ff",x"fb",x"f2",x"c5",x"c0",x"c0",x"ed",x"f6",x"fb",x"ff",x"fa",x"d6",x"d2",x"ce",x"d2",x"db",x"ff",x"ff",x"ff",x"fb",x"f2",x"c4",x"c0",x"c0",x"e9",x"f6",x"ff",x"ff",x"ff",x"fb",x"ed",x"c0",x"e0",x"e0",x"c0",x"f2",x"fb",x"ff",x"ff",x"ff",x"f6",x"cd",x"c4",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"c9",x"cd",x"f2",x"f7",x"ff",x"ff",x"ff",x"fb",x"f6",x"ed",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"c4",x"84",x"48",x"49",x"6d",x"72",x"92",x"96",x"b7",x"b7",x"bb",x"bb",x"db",x"df",x"df",x"df",x"ff",x"ff",x"ff",x"df",x"df",x"df",x"df",x"db",x"db",x"db",x"db",x"d7",x"d7",x"b6",x"92",x"92",x"92",x"6e",x"6e",x"49",x"49",x"25",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"24",x"24",x"24",x"48",x"48",x"49",x"69",x"69",x"49",x"49",x"69",x"6d",x"6d",x"6d",x"6e",x"8e",x"6e",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b7",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b7",x"b6",x"92",x"92",x"6d",x"49",x"24",x"00",x"00",x"00",x"20",x"6e",x"ff",x"db",x"b2",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"b6",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"29",x"24",x"24",x"24",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"a0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c5",x"f2",x"ff",x"ff",x"ff",x"ff",x"d1",x"a4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"ed",x"fb",x"ff",x"ff",x"ff",x"d2",x"a9",x"84",x"a4",x"c5",x"c9",x"ed",x"e9",x"c4",x"a0",x"a0",x"ed",x"f7",x"ff",x"ff",x"ff",x"fa",x"ad",x"a9",x"c9",x"c9",x"c4",x"c4",x"a4",x"a8",x"d1",x"fa",x"ff",x"ff",x"ff",x"f6",x"c4",x"c0",x"c5",x"f6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f2",x"e9",x"c0",x"c0",x"c4",x"ed",x"f6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"f6",x"e9",x"c0",x"c0",x"c0",x"e9",x"f2",x"ff",x"ff",x"ff",x"f6",x"e9",x"e0",x"e0",x"e0",x"c0",x"c9",x"f2",x"ff",x"ff",x"ff",x"ff",x"da",x"d1",x"c8",x"c4",x"c0",x"c0",x"a0",x"a0",x"c4",x"c4",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c4",x"ed",x"f6",x"ff",x"ff",x"ff",x"ff",x"d6",x"c9",x"c0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c4",x"84",x"69",x"6d",x"72",x"72",x"92",x"96",x"97",x"b7",x"97",x"b7",x"b7",x"bb",x"db",x"db",x"d7",x"d7",x"b7",x"b6",x"92",x"92",x"72",x"6e",x"6e",x"69",x"49",x"49",x"25",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b7",x"b6",x"92",x"92",x"6d",x"49",x"24",x"00",x"00",x"00",x"00",x"69",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"da",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"29",x"24",x"24",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"a0",x"e0",x"e0",x"e0",x"e0",x"c0",x"e5",x"f2",x"ff",x"ff",x"ff",x"ff",x"f2",x"c9",x"c0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"e4",x"e4",x"e4",x"e0",x"e0",x"c0",x"e9",x"fb",x"ff",x"ff",x"ff",x"f7",x"f2",x"d1",x"f2",x"f6",x"f6",x"f6",x"f2",x"e9",x"c0",x"a4",x"f2",x"fb",x"ff",x"ff",x"fb",x"f2",x"c4",x"c0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"e9",x"f6",x"fb",x"ff",x"ff",x"f6",x"c8",x"a4",x"c4",x"f2",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fa",x"f6",x"ed",x"e4",x"c0",x"c0",x"c4",x"e9",x"f6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f2",x"c4",x"c0",x"c0",x"c0",x"c5",x"f2",x"ff",x"ff",x"ff",x"f6",x"c9",x"c0",x"e0",x"e0",x"c0",x"c4",x"ed",x"f6",x"ff",x"ff",x"ff",x"ff",x"f6",x"f2",x"ed",x"c9",x"c9",x"c9",x"cd",x"d1",x"cd",x"e9",x"e4",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c4",x"c9",x"f6",x"ff",x"ff",x"ff",x"fb",x"ce",x"c4",x"e0",x"e0",x"e0",x"e0",x"e4",x"c4",x"84",x"64",x"49",x"4d",x"4d",x"49",x"4d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"45",x"45",x"25",x"25",x"24",x"24",x"24",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"28",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b7",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"24",x"00",x"00",x"00",x"25",x"b6",x"db",x"ff",x"ff",x"ff",x"db",x"b7",x"6e",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"40",x"a0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e5",x"f2",x"fb",x"ff",x"ff",x"ff",x"f6",x"ed",x"c4",x"c0",x"c0",x"c0",x"c0",x"c4",x"c9",x"ed",x"f2",x"ed",x"e9",x"c0",x"c0",x"c9",x"fb",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"fa",x"e9",x"c4",x"c5",x"f2",x"fb",x"ff",x"ff",x"f6",x"e9",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"e4",x"ed",x"f6",x"fb",x"fa",x"f1",x"c4",x"a4",x"c4",x"ed",x"f2",x"f6",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"f6",x"f1",x"c9",x"e4",x"e0",x"e0",x"e0",x"c0",x"e4",x"ed",x"f2",x"f6",x"fb",x"ff",x"ff",x"ff",x"ff",x"fb",x"fa",x"f6",x"f2",x"e9",x"c0",x"c0",x"c0",x"c0",x"c4",x"ed",x"fa",x"ff",x"ff",x"f6",x"c9",x"c0",x"e0",x"e0",x"e0",x"e0",x"e9",x"f2",x"f7",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"d6",x"f6",x"f6",x"f6",x"fb",x"fa",x"f2",x"e5",x"e0",x"c0",x"a0",x"a4",x"a4",x"c4",x"c4",x"c0",x"c0",x"c0",x"a0",x"ee",x"fb",x"ff",x"ff",x"fb",x"f2",x"e5",x"e0",x"e0",x"e0",x"e0",x"e4",x"c0",x"80",x"40",x"24",x"24",x"24",x"24",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"24",x"00",x"00",x"00",x"00",x"25",x"69",x"92",x"ff",x"ff",x"b7",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"6d",x"69",x"49",x"49",x"49",x"24",x"24",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"40",x"20",x"40",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"ee",x"fb",x"ff",x"ff",x"ff",x"fb",x"f6",x"ce",x"c9",x"a5",x"a9",x"a9",x"ad",x"d2",x"fa",x"fb",x"fb",x"f2",x"c4",x"a0",x"cd",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fa",x"e9",x"e4",x"e5",x"f2",x"fb",x"ff",x"fb",x"f2",x"e5",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"ed",x"ee",x"ed",x"e9",x"c4",x"c0",x"c0",x"e4",x"e5",x"e9",x"ed",x"ed",x"ed",x"ed",x"e9",x"e9",x"e9",x"e4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e9",x"ed",x"f2",x"f6",x"f6",x"f2",x"f2",x"ed",x"e5",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e5",x"ee",x"f2",x"f2",x"ed",x"e4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e5",x"ee",x"f6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"f6",x"e9",x"e0",x"c0",x"c8",x"f2",x"f7",x"f6",x"cd",x"c4",x"a0",x"a0",x"80",x"cd",x"fa",x"ff",x"ff",x"ff",x"f2",x"e5",x"c0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"40",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"28",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b7",x"b6",x"b6",x"92",x"71",x"6d",x"49",x"25",x"24",x"00",x"00",x"00",x"00",x"20",x"25",x"6e",x"6e",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"6d",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"69",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"40",x"40",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"60",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c9",x"f2",x"fb",x"ff",x"ff",x"ff",x"fb",x"fb",x"d6",x"d6",x"d6",x"d6",x"db",x"ff",x"ff",x"ff",x"fb",x"f2",x"a4",x"a0",x"c9",x"f6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"da",x"f6",x"f2",x"e9",x"e0",x"c0",x"e9",x"ed",x"d1",x"cd",x"c9",x"e4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c4",x"c4",x"c4",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"c4",x"c4",x"c4",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e9",x"e9",x"c4",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c4",x"ed",x"f2",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f2",x"e4",x"c0",x"c0",x"ed",x"f6",x"ff",x"ff",x"f6",x"f1",x"ed",x"cd",x"cd",x"f6",x"fb",x"ff",x"ff",x"ff",x"f2",x"e5",x"c0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"40",x"20",x"40",x"40",x"60",x"60",x"40",x"40",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"40",x"40",x"60",x"80",x"a0",x"a0",x"a0",x"80",x"60",x"60",x"40",x"40",x"60",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c4",x"cd",x"f6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"f6",x"cd",x"a4",x"a0",x"c9",x"f2",x"f6",x"f6",x"f6",x"f6",x"f6",x"d6",x"f2",x"ed",x"cd",x"cd",x"c9",x"e0",x"e0",x"e0",x"c0",x"c4",x"c4",x"c4",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"e0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c4",x"c9",x"d2",x"f6",x"f6",x"fb",x"ff",x"ff",x"fb",x"fb",x"fb",x"f2",x"ed",x"e0",x"c0",x"c0",x"ed",x"f6",x"ff",x"ff",x"ff",x"fb",x"fb",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"fb",x"f2",x"e5",x"c0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"40",x"40",x"60",x"80",x"80",x"a0",x"a0",x"80",x"60",x"60",x"40",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"20",x"20",x"40",x"60",x"80",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"a0",x"80",x"60",x"40",x"40",x"80",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c9",x"f2",x"f6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"f6",x"cd",x"c4",x"c0",x"c0",x"e4",x"e8",x"e8",x"e9",x"c4",x"c4",x"a4",x"a4",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c4",x"c9",x"ed",x"ed",x"ed",x"f2",x"f2",x"f2",x"ed",x"e5",x"e0",x"e0",x"e0",x"c0",x"e5",x"ed",x"f6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"ed",x"e4",x"c0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"40",x"40",x"60",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"84",x"60",x"40",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"04",x"24",x"24",x"24",x"49",x"29",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"48",x"49",x"49",x"49",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"25",x"24",x"00",x"00",x"40",x"60",x"80",x"a0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"60",x"60",x"40",x"80",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c4",x"e9",x"ed",x"f6",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"f2",x"ee",x"e9",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e4",x"c4",x"c0",x"c0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c4",x"c4",x"c0",x"c0",x"c0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"e0",x"e4",x"e4",x"e4",x"e4",x"c4",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c5",x"cd",x"f6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"e9",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"80",x"40",x"40",x"60",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"80",x"80",x"40",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"91",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"72",x"6d",x"49",x"49",x"24",x"00",x"20",x"44",x"84",x"a4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a0",x"80",x"60",x"60",x"60",x"60",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c4",x"e9",x"ee",x"f2",x"f6",x"f6",x"f6",x"f6",x"f2",x"ed",x"e9",x"c5",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a4",x"a4",x"84",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"a4",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a4",x"a4",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"c4",x"c4",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c4",x"ed",x"f2",x"f6",x"fb",x"fb",x"fb",x"fb",x"fb",x"f6",x"f1",x"e9",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"80",x"40",x"40",x"60",x"80",x"a0",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"80",x"44",x"20",x"00",x"00",x"00",x"24",x"24",x"45",x"49",x"49",x"4d",x"6d",x"6d",x"6d",x"91",x"92",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"49",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"69",x"49",x"24",x"00",x"00",x"44",x"84",x"a4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"60",x"60",x"40",x"60",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c4",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"20",x"20",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"84",x"84",x"84",x"84",x"a0",x"a0",x"a4",x"a4",x"a0",x"a0",x"c0",x"c0",x"e4",x"e0",x"e0",x"c0",x"e0",x"e0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c4",x"a4",x"c9",x"e9",x"ed",x"ed",x"e9",x"e5",x"c4",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"40",x"40",x"60",x"80",x"a0",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"80",x"40",x"20",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"6d",x"6d",x"71",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"4d",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"8e",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"96",x"92",x"6d",x"49",x"49",x"24",x"00",x"00",x"20",x"60",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"80",x"60",x"40",x"40",x"60",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"20",x"20",x"20",x"00",x"00",x"20",x"20",x"20",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"00",x"00",x"20",x"20",x"20",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"c4",x"c0",x"c0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"c0",x"e0",x"e0",x"e4",x"e0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"40",x"40",x"60",x"80",x"a0",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"60",x"20",x"20",x"00",x"00",x"24",x"28",x"49",x"49",x"6d",x"6d",x"71",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b7",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b7",x"b6",x"b6",x"92",x"92",x"92",x"91",x"6d",x"71",x"71",x"6d",x"6d",x"6d",x"6d",x"8e",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"6d",x"49",x"49",x"24",x"00",x"00",x"20",x"40",x"80",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"40",x"40",x"40",x"60",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c4",x"c4",x"c4",x"a4",x"a4",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"a0",x"a0",x"c0",x"c0",x"c4",x"c4",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e4",x"e4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"60",x"40",x"40",x"60",x"80",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"40",x"20",x"00",x"00",x"24",x"24",x"49",x"49",x"6d",x"6d",x"91",x"92",x"96",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"6d",x"6d",x"49",x"24",x"20",x"00",x"00",x"00",x"20",x"40",x"80",x"c0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"60",x"40",x"40",x"80",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c4",x"c4",x"c4",x"a4",x"a4",x"a4",x"80",x"60",x"60",x"40",x"40",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"40",x"40",x"40",x"60",x"60",x"80",x"a0",x"a0",x"c4",x"c4",x"a4",x"c4",x"c4",x"c4",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"80",x"40",x"40",x"60",x"80",x"a0",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"c0",x"80",x"40",x"20",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b2",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"92",x"92",x"6d",x"49",x"45",x"24",x"00",x"00",x"00",x"00",x"00",x"60",x"a0",x"c0",x"c0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"60",x"40",x"60",x"80",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"84",x"84",x"64",x"60",x"60",x"40",x"40",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"04",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"80",x"60",x"40",x"60",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"80",x"40",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"6d",x"6e",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"92",x"92",x"6d",x"49",x"49",x"24",x"20",x"00",x"00",x"00",x"00",x"20",x"60",x"80",x"a0",x"c0",x"c0",x"c0",x"c0",x"a0",x"80",x"60",x"60",x"60",x"60",x"a4",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c4",x"c4",x"a0",x"80",x"80",x"80",x"60",x"60",x"40",x"40",x"20",x"20",x"20",x"00",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"a0",x"a0",x"c4",x"c4",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"60",x"60",x"60",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"80",x"60",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"92",x"92",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"40",x"80",x"a0",x"c0",x"c0",x"c0",x"a0",x"80",x"60",x"60",x"60",x"60",x"a4",x"c4",x"c4",x"c0",x"a0",x"a4",x"80",x"80",x"60",x"60",x"40",x"40",x"40",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"40",x"40",x"60",x"60",x"60",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c4",x"a0",x"80",x"60",x"60",x"60",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"80",x"60",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"6d",x"49",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"60",x"a0",x"c0",x"c0",x"c0",x"a0",x"80",x"60",x"60",x"40",x"60",x"84",x"84",x"80",x"80",x"80",x"60",x"40",x"40",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"24",x"24",x"24",x"28",x"28",x"29",x"29",x"49",x"45",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"04",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"60",x"60",x"60",x"60",x"80",x"a0",x"a4",x"80",x"60",x"40",x"40",x"60",x"80",x"80",x"a0",x"c0",x"c0",x"a0",x"60",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"6d",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"60",x"80",x"c0",x"c0",x"a0",x"a0",x"80",x"60",x"60",x"40",x"20",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"04",x"24",x"24",x"24",x"24",x"24",x"28",x"28",x"29",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"29",x"24",x"24",x"24",x"24",x"04",x"04",x"04",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"40",x"40",x"60",x"40",x"40",x"20",x"40",x"60",x"60",x"80",x"a0",x"c0",x"c0",x"a0",x"60",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"6d",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"60",x"a0",x"c0",x"c0",x"a0",x"a0",x"80",x"60",x"40",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"44",x"44",x"44",x"44",x"49",x"49",x"49",x"49",x"49",x"4d",x"4d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"69",x"69",x"69",x"69",x"49",x"49",x"49",x"49",x"49",x"44",x"44",x"24",x"29",x"24",x"24",x"24",x"24",x"24",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"40",x"60",x"80",x"a0",x"c0",x"c0",x"c0",x"a0",x"60",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"6d",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"20",x"40",x"80",x"a0",x"c0",x"c0",x"a0",x"a0",x"80",x"60",x"40",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"49",x"49",x"49",x"69",x"69",x"69",x"69",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"72",x"72",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"69",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"04",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"40",x"60",x"80",x"a0",x"c0",x"e0",x"e0",x"c0",x"80",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"6d",x"6d",x"92",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"6d",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"20",x"40",x"60",x"a0",x"c0",x"c0",x"c0",x"c0",x"a0",x"80",x"60",x"40",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"29",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"8d",x"8d",x"8e",x"8e",x"92",x"92",x"92",x"92",x"92",x"96",x"96",x"96",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"72",x"72",x"72",x"6e",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"40",x"60",x"80",x"a0",x"a0",x"c0",x"e0",x"e0",x"c0",x"a0",x"60",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"96",x"92",x"6d",x"6d",x"49",x"49",x"24",x"20",x"00",x"00",x"00",x"40",x"60",x"a0",x"c0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"60",x"40",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"49",x"49",x"49",x"49",x"4d",x"4d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"b2",x"b2",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"96",x"96",x"96",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"8e",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"40",x"40",x"60",x"a0",x"a0",x"c0",x"c0",x"e0",x"e0",x"c0",x"80",x"40",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"44",x"24",x"00",x"00",x"00",x"00",x"60",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"40",x"40",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"4d",x"4d",x"6d",x"6d",x"6d",x"71",x"71",x"92",x"92",x"92",x"92",x"92",x"92",x"96",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"96",x"96",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"44",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"40",x"60",x"80",x"a0",x"a0",x"c0",x"c0",x"e0",x"e0",x"c0",x"80",x"40",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"92",x"92",x"6d",x"6d",x"49",x"44",x"20",x"00",x"00",x"00",x"20",x"80",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"60",x"40",x"20",x"00",x"00",x"00",x"04",x"04",x"24",x"44",x"49",x"49",x"4d",x"6d",x"6d",x"6d",x"8d",x"92",x"92",x"92",x"92",x"92",x"b2",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b7",x"bb",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"d6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"96",x"92",x"92",x"92",x"92",x"92",x"72",x"6e",x"6d",x"6d",x"4d",x"49",x"45",x"24",x"24",x"04",x"00",x"00",x"00",x"00",x"00",x"20",x"40",x"60",x"80",x"a0",x"a0",x"c0",x"c0",x"e0",x"e0",x"c0",x"a0",x"60",x"20",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"ba",x"96",x"92",x"92",x"6d",x"6d",x"49",x"24",x"00",x"00",x"00",x"20",x"40",x"a0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"60",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"bb",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b7",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"96",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"29",x"24",x"24",x"00",x"00",x"00",x"00",x"20",x"40",x"40",x"60",x"80",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"40",x"00",x"00",x"00",x"00",x"24",x"29",x"49",x"6d",x"8e",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"ba",x"96",x"92",x"8d",x"8d",x"69",x"49",x"04",x"00",x"00",x"20",x"40",x"80",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"60",x"40",x"20",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"ba",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"d6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"8d",x"6d",x"6d",x"49",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"20",x"20",x"40",x"60",x"80",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"60",x"20",x"00",x"00",x"00",x"04",x"24",x"49",x"6d",x"8e",x"92",x"b2",x"b6",x"bb",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"92",x"8d",x"6d",x"49",x"49",x"04",x"00",x"00",x"20",x"60",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a0",x"60",x"40",x"20",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"20",x"20",x"60",x"80",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"60",x"20",x"00",x"00",x"00",x"24",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"da",x"b6",x"92",x"8d",x"6d",x"49",x"29",x"00",x"00",x"20",x"60",x"80",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"60",x"40",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"40",x"60",x"a0",x"c0",x"c0",x"c0",x"c0",x"e0",x"c0",x"c0",x"a0",x"40",x"00",x"00",x"00",x"24",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"bb",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"49",x"28",x"00",x"00",x"40",x"80",x"a0",x"c5",x"c4",x"a0",x"a0",x"80",x"60",x"40",x"40",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"8e",x"6d",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"60",x"60",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"a0",x"60",x"20",x"00",x"00",x"24",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"49",x"24",x"00",x"00",x"40",x"84",x"a0",x"a0",x"60",x"40",x"40",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b2",x"92",x"92",x"6d",x"6d",x"49",x"49",x"28",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"40",x"40",x"60",x"80",x"a4",x"a4",x"84",x"40",x"00",x"00",x"24",x"49",x"6d",x"71",x"92",x"b6",x"b6",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"96",x"92",x"6d",x"49",x"24",x"00",x"00",x"40",x"60",x"60",x"60",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"45",x"49",x"49",x"49",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"4d",x"49",x"49",x"24",x"24",x"24",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"40",x"60",x"60",x"60",x"40",x"00",x"00",x"24",x"49",x"6d",x"71",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"ba",x"b6",x"96",x"92",x"8d",x"69",x"44",x"00",x"00",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"45",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"d6",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"6d",x"4d",x"49",x"49",x"24",x"24",x"24",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"00",x"00",x"24",x"4d",x"6d",x"92",x"96",x"b6",x"b6",x"db",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"8e",x"6d",x"69",x"24",x"20",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"04",x"24",x"24",x"24",x"29",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"48",x"44",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"49",x"6d",x"72",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"49",x"44",x"24",x"24",x"04",x"04",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"4d",x"4d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"69",x"69",x"49",x"48",x"24",x"24",x"24",x"24",x"04",x"04",x"00",x"00",x"20",x"20",x"20",x"24",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"49",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"4d",x"6d",x"6d",x"6d",x"71",x"91",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"72",x"6d",x"8d",x"6d",x"6d",x"49",x"49",x"45",x"45",x"45",x"29",x"29",x"25",x"24",x"24",x"44",x"49",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"d7",x"b6",x"96",x"92",x"72",x"71",x"6d",x"6d",x"6d",x"6d",x"49",x"4d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"91",x"92",x"92",x"91",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"6d",x"4d",x"4d",x"6d",x"69",x"69",x"69",x"4d",x"4d",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"92",x"b2",x"b6",x"b6",x"d7",x"db",x"df",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"db",x"db",x"b6",x"b6",x"96",x"92",x"92",x"92",x"91",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6e",x"92",x"92",x"92",x"92",x"b2",x"b2",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"db",x"db",x"db",x"d6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"72",x"72",x"71",x"8d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"72",x"72",x"92",x"92",x"b6",x"b6",x"d6",x"db",x"db",x"df",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff")
);

constant object : object_form := (
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000011111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000001111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000011111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111110011111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111110011111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000001111111111111111111111111111111111000000000000001111111111111111111111111111111111100011111111111111111111000000000000000000000000000000111111111111111111000000000000000000000000001111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000011111111111111111111100000000000000000000000000000000000000000000000111111111111111111111111111111111111100000000000011111111111111111111111111111111111000001111111111111111111110000000000000000000000011111111111111111111111111110000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000001111111111111111111111111111111111111111100000000111111111111111111111111111111111111000001111111111111111111111100000000000000000111111111111111111111111111111111111110000011111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000011111111111111111111111111111111111111111111111111001111111111111111111111111111111111110000001111111111111111111111110010000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000111111111111111111111111111111000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000111111111111111111111111111000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000011111111111111111111111111111111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111111111111111111111111000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000011111111111111111111111111111111111111111111110000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111100100000000111000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111110111111111111111111111111000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000111111111111111001111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111111111111111100011111111111111111111111110000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000111111111111111101111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000001111111111111111100111111111100111111111111101111111111111110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111111111111111111000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000111111111111111110111111111111111111111111111111111111111111111100011111111111111111111110000000000011111111111111111111111111111111111111111111111111111111000001111111111111111111111111100000000000000000011111111111111111111110011111111111111111001111111111111111111111111111111111110000000000000000000000000000000000000000111111111111111111111111111111111000011111111111111111111111111111111111111111111000111111111111111111111111111111000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111111111111111111110000000000000000111111111111111110001111111111111111111111000111111111111111111111111111111111111100000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111100011111111111111011111111111111111111111100000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111110000011111111111111111111111111110000000000000000111111111111111110011111111111111111111111000111111111111111111111111111111111111110000000000000000000000000000000000001111111111111111111111111110011111111111111111111111111111111111111111110011111111111111111110011111111111111111111100000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000111111111111111111100011111111111111111111111111111111111111111111111111101111111111111111111111111111111111101111111111111111111111111111111111111111001100000010001111111111111111111111111000000000000001111111111111111100111111111111111111111111001111111111111111111111111111111111111111000000000000000000000000000000000111111111111111111111111111001111111111111111111111111011111111111111110011111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000001111111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111110000000000001111111111111111101111111111111111111111111011111111111111111111111111111111111111111100000000000000000000000000000011111111111111111111111111000111111111111111111111111111110111111111111011111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000011111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000011111111111111111111110000000000011111111111111111101111111111111111111111110011111111111111111111111111111111111111111110000000000000000000000000000111111111111111111111111110011111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000011111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111100000000000000000001111111111111111111111111000000000011111111111111111011111111111111111111111110011111111111111111111111111111111111111111110000000000000000000000000011111111111111111111111111101111111111111111111111111111111111111111111001111111111111111111111111111111111011111111111111110000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000111111111111111111111111111111111111100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111110000000000001000011111111111111111111111111000000000011111111111111111011111111111111111111111100111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111111110011111111111111111111111111111111111101111110111111111111111111111111111111111111011111111111111110000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000011111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111000000000000000111111111111111111111111111100000000111111111111111110111111111111111111111111100111111111111111111111111111111111111111111110000000000000000000000011111111111111111111111111100111111111111111111111111111111111111110111101111111111111111111111111111111111111101111111111111110000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000001111111111111111111111111111111111111111111111000000000011111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111100000000000001111111111111111111111111111100000000111111111111111110111111111111111111111111001111111111111111111111111111111111111111111100000000000000000000000111111111111111111111111111001111111111111111111111111111111111111110111111111111111111111111111111111111111111101111111111111110000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000011111111111111111111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111100000000000001111111111111111111111111111110000001111111111111111100111111111111111111111111011111111111111111111111111111111111111111111100000000000000000000000111111111111111111111111111011111111111111111111111111111111111111110001111111111111111111111111111111111111111100111111111111110000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111000001111111111111111111111111111111111100001111111111111111111111111111110111111111111111111111111111111111100000000000001111111111111111111111111111111011111111111111111111101111111111111111111111110011111111111111111111111111111111111111111111100000000000000000000000111111111111111111111111110111111111111111111111111111111111111111110011111111111111111111111111111111111111111101111111111111110000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111110000111111111111111111111111111111100000000011111111111111111111111111100111111111111111111111111111111111100000000000001111111111111111111111111111111111111111111111111111001111111111111111111111110011111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111101111111111111111111111111111111111111111100011111111111111111111111111111111111111111101111111111111110000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111000111111001111111111111111111111111100111111111111111111111111111111111000000000000011111111111111111111111111111111111111111111111111111011111111111111111111111110111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111011111111111111111111111110011111111111111100111111111111111111111111100111111111111111001111111111111110000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111110011111111101111111111111111111111111100111111111111111111111111111111111000011111000011111111111111111111111111111111111111111111111111110011111111111111111111111100111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111110011111111111111111111111100011111111111111100111111111111111111111111000011111111111111001111111111111110000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111100111111111111111111111111111111111111101111111111100011111111111111111111011111111110001111111111111111111111111111111111111111111111111110111111111111111111111111101111111111111111111111111111111111111111111111000000000000111000000000011111111111111111111110111111111111111111111111100111111111111111001111111111111111111111111000111111111111111011111111111111110000000000000001111111100000000000000000000000000000000"),
("0000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111001111111111100111111111111111111111111001111111111111111111111111111111110011111111111100111111111111111111111111111111111111111111111111100111111111111111111111111001111111111111111111111111111111111111111111111000000001111111000000000011111111111111111111100111111111111111111111111000111111111111111001111111111111111111111110001111111111111110011111111111111110000000001111111111111111110000000000000000000000000000"),
("0000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111001111111111101111111111111111111111111001111110111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111101111111111111111111111111011111111111111111111111111111111111111111111110000001111111111100100000011111111111111111111101111111111111111111111110000111111111111110011111111111111111111111110001111111111111110111111111111111111110001111111111111111111111000000000000000000000000000"),
("0000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111110011111111111101111111111111111111111110011110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111110011111111111111111111111111111111111111111111110000111111111111111100000001111111111111111111001111111111111111111111110001111111111111110111111111111111111111111110011111111111111100111111111111111111111111111111111111111111111100000000000000000000000000"),
("0000000000000000011111111111111111111111110011111111111111111111111111111111111111111111111111110111111111111111111111111110111111111111001111111111111111111111110111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111100111111111111111111110000001111111111111111111011111111111111111111111110001111111111111100111111111111111111111111100011111111111111101111111111111111111111111111111111111111111111111000000000000000000000000"),
("0000000000000000111111111111111111111111110111111111111111111111111111111111111111111111111111100111111111111111111111111100111111111111011111111111111111111111110011011111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111011111111111111111111111110001111111111111111110011111111111111111111111100011111111111111101111111111111111111111111100011111111111111001111111111111111111111111111111111111111111111111110000000000000000000000"),
("0000000000000001111111111111111111111111100111111111111111111111111111111111111111111111111111101111111111111111111111111101111111111110011111111111111111111111100100111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111000111111111111111110111111111111111111111111000111111111111111001111111111111111111111111000111111111111111001111111111111111111111111111111111111111111111111111000000000000000000000"),
("0000000000000111111111111111111111111111000011111111111111111111111111111111111111111111111111001111111111111111111111111001111111111110111111111111111111111111000001111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111101111111111111111111111111000111111111111111001111111111111111111111111001111111111111110011111111111111111111111111111111111111111111111111111110000000000000000000"),
("0000000000001111111111111111111111111111000011111111111111111111111111111111111111111111111111011111111111111111111111110011111111111101111111111111111111111111000001111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111001111111111111110011111111111111111111111110001111111111111110011111111111111111111111111111111111111111111111111111111000000000000000000"),
("0000000000001111111111111111111111111110000001111111111111111111111111111111111111111111111110111111111111111111111111110011111111111101111111111111111111111111000011111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111001111111111111111111111110001111111111111110011111111111111111111111110001111111111111100111111111111111111111111111111111111111111111111111111111110000000000000000"),
("0000000000011111111111111111111111111110000001111111111111111111111111111111111111111111111110111111111111111111111111110011111111111001111111111111111111111110000011111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111110001111111111111110011111111111111111111111100011111111111111100111111111111111111111111111111111111111111111111111111111110000000000000000"),
("0000000001111111111111111111111111111000000000111111111111111111111111111111111111111111111101111111111111111111111111100111111111111011111111111111111111111110100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111110011111111111111100111111111111111111111111100011111111111111101111111111111111111111111111111111111111111111111111111111111110000000000000"),
("0000000001111111111111111111111111111000000000111111111111111111111111111111111111111111111101111111111111111111111111101111111111111011111111111111111111111100110011111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111100011111111111111100111111111111111111111111000111111111111111001111111111111111111111111111111111111111111111111111111111111111000000000000"),
("0000000001111111111111111111111111110000000000111111111111111111111111111111111111111111111111111111111111111111111111001111111111110111111111111111111111111100111011111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111100111111111111111001111111111111111111111111000111111111111111011111111111111111111111111111111111111111111111111111111111111111100000000000"),
("0000000011111111111111111111111111110000000000111111111111111111111111111111111111111111111011111111111111111111111111001111111111100111111111111111111111111001111011111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111000111111111111111001111111111111111111111110001111111111111110011111111111111111111111111111111111111111111111111111111111111111110000000000"),
("0000000011111111111111111111111111100000000000011111111111111111111111111111111111111111111011111111111111111111111111011111111111101111111111111111111111111011111001111111111111111111100001111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111110001111111111111110011111111111111111111111110001111111111111100111111111111111111111111111111111111111111110011111111111111111111110000000000"),
("0000000011111111111111111110000000000000000000000000000000110111111111111111111111111111110111111111111111111111111111111111111111101111111111111111111111110011111100111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111110001111111111111110011111111111111111111111100011111111111111100111111111111111111111111111111111111111111110011111111111111111111111000000000"),
("0000000011111111111100000000000000000000000000000000000000011111111111111111111111111111110111111111111111111111111100111111111111011111111111111111111111110011111111000111111111100000011111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111110011111111111111100111111111111111111111111100011111111111111101111111111111111111111111111111111111111111110001111111111111111111111000000000"),
("0000000011111111111110000000000000000000000000000000000000111111111111111111111111111111101111111111111111111111111100111111111111011111111111111111111111100111111111100000000000000001111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111100011111111111111100111111111111111111111111000111111111111111001111111111111111111111111111111111111111111110000111111111111111111111100000000"),
("0000000011111111111111000000000000000000000000000000000001111111111111111111111111111111101111111111111111111111111101111111111110111111111111111111111111101111111111111000000000011111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111000111111111111111001111111111111111111111111000111111111111111011111111111111111111111111111111111111111111110000111111111111111111111100000000"),
("0000000011111111111111100000000000000000000000000000000011111111111111111111111111111111011111111111111111111111111011111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111000111111111111111011111111111111111111111110001111111111111110011111111111111111111111111111111111111111111110000011101110111111111111100000000"),
("0000000011111111111111111000000000000000000000000000001111111111111111111111111111111111011111111111111111111111111011111111111101111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111001111111111111110011111111111111111111111110001111111111111110011111111111111111111111111111111111110010000000000000000000011111111111100000000"),
("0000000011111111111111111000000000000000000000000000011111111111111111111111111111111110011111111111111111111111110011111111111101111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111110001111111111111110111111111111111111111111110011111111111111100111111111111111111111111111111111111111000000000000000000000111111111111100000000"),
("0000000001111111111111111110000000000000000000000001111111111111111111111111111111111110111111111111111111111111110111111111111001111111111111111111111110011110111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111011111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111100011111111111111100111111111111111111111111100111111111111111101111111111111111111111111111111111111111110000000000000000011111111111111100000000"),
("0000000001111111111111111111000000000000000000000011111111111111111111111111111111111101111111111111111111111111100111111111111011111111111111111111111100111100001111111111111111111111111111000011111111111111111111111111111111111111111111111111111111110011111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111100011111111111111100111111111111111111111111000111111111111111101111111111111111111111111111111111111111111100000000000000111111111111111100000000"),
("0000000001111111111111111111000000000000000000000111111111111111111111111111111111111111111111111111111111111111100111111111110011111111111111111111111100111011111111111111111111111111111111011111111111111111111111111000011100100011111111111111111111110111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111100111111111111111001111111111111111111111111001111111111111110111111111111111111111111111111111111111111111110000000010001111111111111111100000000"),
("0000000000111111111111111111000000000000000000000111111111111111111111111111111111111011111111111111111111111111001111111111110111111111111111111111111001111011111111111111111111111111111110111111111111111111111110111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111000111111111111110001111111111111111111111110011111111111111110011111111111111111111111111111111111111111111111110000000001111111111111111100000000"),
("0000000000111111111111111111000000000000000000001111111111111111111111111111111111111011111111111111111111111111001111111111100111111111111111111111111001111111111111011111111111111111111110111111111111111111111111111111111111111111111111111111111111101111111111111111111111111000011111111111111111111111111111111111111111111111111111110111111111111111111111111111111111101111111111111111111111111001111111111111110001111111111111111111111110011111111111111100111111111111111111111111111111111111111111111111100000000001111111111111111100000000"),
("0000000000111111111111111111000000000000000000001111111111111111111111111111111111110011111111111111111111111110011111111111101111111111111111111111111011110111111111111111111111111111111100111111111110111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111110001111111001111111111111111111111110011111111111111100011111111111111111111111110111111111111111101111111111111111111111111111111111111111111111111100010000000111111111111111100000000"),
("0000000000011111111111111110000000000000000000000111111111111111111111111111111111110111111111111111111111111110011111111111101111111111111111111111110011110111111111111111111111111111111101111111111111111111111111111111111111111111110111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111011111111111111111111111111111111111111111100111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111100000000000011111111111111100000000"),
("0000000000111111111111111110000000000000000000000111111111111111111111111111111111100111111111111111111111111100111111111111011111111111111111111111110111101111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111011111111111111111111111110111111111111111111111111011111111111111110011111110011111111111111111111111111111111111111111000111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111100000111100011111111111111100000000"),
("0000000000111111111111111110000000000000000000000111111111111111111111111111111111101111111111111111111111111100111111111110011111111111111111111111100111001111111111111111111111111111111011111111111111111111111111111111111111111111111011111111111110011111111111111111111111111111111111111111101111111111111111111111001111111111111111111111111110111111111111110011111110111111111111111111111111111111111111111110001111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111100011111111001111111111111100000000"),
("0000000000111111111111111100000000011100000000000111111111111111111111111111111111011111111111111111111111111001111111111110111111111111111111111111101111011111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111110111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111100001111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111000111111111101111111111111100000000"),
("0000000000111111111111111000000000111111000000000111111111111111111111111111111111011111111111111111111111111011111111111110111111111111111111111111001111011111111111111111111110011111111111111111111111111111111111111111111111111111111001111111111101111111111111111111111111111111111111111111110111111111111111111101111111111111111111111111111111111111111111100111111101111111111111111111111111111111111111111000011111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111001111111111111111111111111100000000"),
("0000000001111111111111111000000001111111110000000111111111111111111111111111111111111111111111111111111111110011111111111101111111111111111111111111011111111111111111111111111110011111101111111111111111111111111111111111111111111111111101111111111101111111111111111111111111111111111111111111111011111111111111110011111111111111111111111111111111111111111111101111111101111111111111111111111111111111111111110000111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111100000000"),
("0000000001111111111111111000001111111111111000000111111111111111111111111111111110111111111111111111111111110011111111111101111111111111111111111110011111111111111111111111111110011111101111111111111111111111111111111111111111111111111101111111111001111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111001111111011111111111111111111111111111111111111100000111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000"),
("0000000001111111111111111000111111111111111100000111111111111111111111111111111100111111111111111111111111110111111111111011111111111111111111111110011101111111111111111111111110111111101111111111111111111111111111111111111111111111111101111111111011111111111111111111111111111111111111111111111011111111111111011111111111111111111111111111111111111111111111011111110011111111111111111111111111111111111111000000111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000"),
("0000000001111111111111110011111111111111111111001111111111111111111111111111111101111111111111111111111111100111111111111011111111111111111111111100111101111111111111111111111100111111011111111111111111111111111101111111111111111111111101111111111011111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111110011111110111111111111111111111111111111111111110001101111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000"),
("0000000001111111111111100111111111111111111111100111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111100111011111111111111111111111100111110011111111111111111111111110000111111111111111111111101111111110111111111111111111111111110001111111111111111111011111111111101111111111111111111100011111111111111111111111110111111110111111111111111111111111111111111111100111101111111111111111111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000"),
("0000000001111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111001111111111111111111111111111111111111001111011111111111111111111111001111110111111111111111111111111100000111111111111111111111101111111101111111111111111111111111100001111111111111111111011111111111011111111111111111111000001111111111111111111111100111111101111111111111111111111111111111111111001111101111111111111111111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000"),
("0000000000111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111011111111111101111111111111111111111111001110111111111111111111111111011111110111111111111111111111111100001111111111111111111111101111111101111111111111111111111111000001111111111111111111011111111110111111111111111111110011011111111111111111111111000111111101111111111111111111111111111111111100011111011111111111111111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000"),
("0000000000111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111110011111111111101111111111111111111111110011110111111111111111111111110011111101111111111111111111111111000011111111111111111111111001111111101111111111111111111111110010011111111111111111111011111111101111111111111111111110010011111111111111111111111001111111011111111111111111111111111111111111000111111111111111111111111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000"),
("0000000000111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111110111111111111001111111111111111111111100111100111111111111111111111110011111101111111111111111111111111000011111111111111111111111001111111011111111111111111111111110010011111111111111111111011111111111111111111111111111100100011111111111111111111111011111111011111111111111111111111111111111100001111110111111111111111111111111111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000"),
("0000000000111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111100111111111111111111111111111111111111100111101111111111111111111111100111111111111111111111111111111110010111111111111111111111111011111111011111111111111111111111100011111111111111111111110011111110111111111111111111111100111111111111111111111111110011111110111111111111111111111111111111111000111111110111111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000"),
("0000000000111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111101111111111111111111111111111111111111001111011111111111111111111111100111111011111111111111111111111110100111111111111111111111111011111111111111111111111111111111100011111111111111111111110011111110111111111111111111111000011111111111111111111111110011111110111111111111111111111111111111100011111111111111111111111111111111111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000"),
("0000000000111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111001111111111101111111111111111111111110011111011111111111111111111111001111110111111111111111111111111100100111111111111111111111110011111111111111111111111111111111100001111111111111111111110111111101111111111111111111111010011111111111111111111111110111111100111111111111111111111111111110000111111111111111111111111111111111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000"),
("0000000000111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111011111111111111111111111111111111111100011111011111111111111111111111001111110111111111111111111111111100101111111111111111111111110111111101111111111111111111111111000001111111111111111111100111111101111111111111111111111011011111111111111111111111100111111101111111111111111111111111110000011111111111001111111111111111111111111110000111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111000000000000000"),
("0000000000011111111111111111111111111111111111111111111111111111111111111110011111111111111111111111110011111111111111111111111111111111111000111110111111111111111111111110011111111111111111111111111111111000001111111111111111111111100111111101111111111111111111111111000011111111111111111111100111111011111111111111111111110010111111111111111111111111001111111111111111111111111111111111000001111111111111011111111111111111111111111000011111111111111111111111111111111111111111111111111111110111111111111111111111111111111111110000000000000000"),
("0000000000001111111111111111111111111111111111111111111111111111111111111110111111111111111111111111110011111111011111111111111111111111111001111101111111111111111111111110011111101111111111111111111111111000011111111111111111111111100111111001111111111111111111111110010011111111111111111111100111110111111111111111111111110001111111111111111111111111001111111111111111111111111111111110000111111111111110111111111111111111111111100000111111111111111111111111111111111111111100000011111111110111111111111111111111111111111100000000000000000000"),
("0000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111110011111101111111111111111111111110111111101111111111111111111111111000011111111111111111111111001111111011111111111111111111111100010111111111111111111111101111110111111111111111111111101101111111111111111111111111011111110111111111111111111111111100111111111111111110111111111111111111111111100111111111111111111111111111111111111111100000000001111111110111111111111111111111111111111000000000000000000000"),
("0000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111100111111001111111111111111111111100111111011111111111111111111111110000111111111111111111111111001111110111111111111111111111111100111111111111111111111111011111111111111111111111111111101101111111111111111111111110011111110111111111111111111111111100111111111111111100111111111111111111111111101111111111111111111111111111111111111110000111111001111111110111111111111111111111111111100000000000000000000000"),
("0000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111001111111111111111111111111111111100111110011111111111111111111111110000111111111111111111111111011111110111111111111111111111111100101111111111111111111111011111101111111111111111111111001111111111111111111111111110111111110111111111111111111111111101111111111111111101111111111111111111111111001111111111111111111111111111111111110000111111111101111111110111111111111111111111100000000000000000000000000000"),
("0000000000000000011111111111111111111111111111111111111111111111111111111011111111111111111111111111000011111111111111111111111111111110011111111011111111111111111111111001111110111111111111111111111111100001111111111111111111111110011111111111111111111111111111111000101111111111111111111110011111011111111111111111111111011111111111111111111111111100111111111111111111111111111111111001111111111111111001111111111111111111111110011111111111111111111111111111111111100011111111111111111111110111111111111111111100000000000000000000000000000000"),
("0000000000000000001111111111111111111111111111111111111111111111111111111011111111111111111111111111001111111111111111111111111111111000111111111111111111111111111111111001111111111111111111111111111111100001111111111111111111111110111111101111111111111111111111111010011111111111111111111110111111011111111111111111111110011011111111111111111111111101111111111111111111111111111111111011111111111111111011111111111111111111111110011111111111111111111111111111111111000111111111111101111111100111111111111111111000000000000000000000000000000000"),
("0000000000000000000001111111111111111111111111111111111111111111111111110111111111111111111111111110111111111111111111111111111111100001111111111111111111111111111111110011111101111111111111111111111111000011111111111111111111111100111111101111111111111111111111110010111111111111111111111100111110111111111111111111111110010011111111111111111111111101111111011111111111111111111111110011111111111111111111111111111111111111111100111111111111111111111111111111111110011111111111111101111111100111111111111111110000000000000000000000000000000000"),
("0000000000000000000000001111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111110000111111111101111111111111111111111110111111101111111111111111111111111000011111111111111111111111101111111011111111111111111111111110010111111111111111111111001111110111111111111111111111100010111111111111111111111111001111111011111111111111111111111110111111111111111110111111111111111111111111100111111111111111111111111111111111001111111111111111111111111100111111111111111100000000000000000000000000000000000"),
("0000000000000000000000000000111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111100111111011111111111111111111111110000111111111111111111111111001111110111111111111111111111111100001111111111111111111111001111100111111111111111111111100011111111111111111111111110011111110111111111111111111111111100111111111111111100111111111111111111111111001111111111111111111111111111111110001111111111111111111111111101111111111111111000000000000000000000000000000000000"),
("0000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111111111111111111111111111100111111011111111111111111111111110000111111111111111111111111011111110111111111111111111111111100101111111111111111111111001111101111111111111111111111000011111111111111111111111110011111110111111111111111111111111101111111111111111101111111111111111111111111001111111111111111111111111111111100111111111111111111111111111001111111111111111000000000000000000000000000000000000"),
("0000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111111011111111111111111111111001111110111111111111111111111111100001111111111111111111111110011111100111111111111111111111111001101111111111111111111110011111001111111111111111111111001001111111111111111111111100111111101111111111111111111111111001111111111111111111111111111111111111111111011111111111111111111111111111111001111111111111111111111111111001111111111111111000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111000001111111111111110011111111111111111111111001111110111111111111111111111111100001111111111111111111111110011111101111111111111111111111111001101111111111111111111110011111011111111111111111111110011011111111111111111111111100111111101111111111111111111111111001111111111111111011111111111111111111111110011111111111111111111111111111110001111111111111111111111111111011111111111111110000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000011111111111111111111110111111111111111111111111111111111111111111111110000001111111111111111101111111111111111111111110011111101111111111111111111111111100001111111111111111111111100111111111111111111111111111111110010011111111111111111111110111110111111111111111111111110010111111111111111111111111001111111011111111111111111111111110011111111111111111011111111111111111111111110111111111111111111111111111111110011111111111111111111111111111011111111111111110000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000111111111111111111110111111111111111111111111111111111111111111100000001111111111111111111101111111111111111111111110011111101111111111111111111111111000011111111111111111111111100111111011111111111111111111111110010111111111111111111111111111110111111111111111111111100110111111111111111111111111011111111011111111111111111111111110111111111111111110111111111111111111111111100111111111111111111111111111111100111111111111111111111111111110011111111111111110000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111110000000000111111111111111111111111111111111111111111111110111111111111111111111111111111111000011111111111111111111111001111111011111111111111111111111110000111111111111111111111111111111111111111111111111111101111111111111111111111111110011111111111111111111111111111111100111111111111111101111111111111111111111111100111111111111111111111111111111001111111111111111111011111111110111111111111111110000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111111111101111111111111111111111111111111110000111111111111111111111111001111110111111111111111111111111100001111111111111111111111111111111111111111111111111111100001111111111111111111111110011111111111111111111111111111111100111111111111111111111111111111111111111111001111111111111111111111111111110001111111111111111111111111111100111111111111111100000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000011111111111111111011111111111111111111111111000000000001111111111111111111111111111111111111111111111111111111111001111110111111111111111111111111110000111111111111111111111110011111111111111111111111111111111000001111111111111111111111111111111111111111111111111111000011111111111111111111111100111111111111111111111111111111111001111111111111111111111111111111111111111111011111111111111111111111111111100011111111111111111111111111111001111111111111111100000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000011111111111111111011111111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111100001111111111111111111111110111111111111111111111111111111111001111111111111111111111111111111111111111111111111111110010011111111111111111111111101111111111111111111111111111111111011111111111111111111111111111111111111111110011111111111111111111111111111000111111111111111111111111111111011111111111111111000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000011111111111111110011111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111000111111111111111111111111111111100001111111111111111111111110111111111111111111111111111111110011111111111111111111111111111111111111111111111111111110010111111111111111111111111100111111111111111111111111111111111011111111111111111111111111111111111111111110111111111111111111111111111110001111111111111111111111111111110011111111111111111000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000111111111111111110111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111000011111111111111111111111111011111111111111111111111111111110010111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111110011111111111111111111111111100011111111111111111111111111111100111111111111111110000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111100111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111000011111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111111111111111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111000111111111111111111111111111111100111111111111111100000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111111111111111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111111111111111111111111001111111111111111100000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110010111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111110011111111111111111100000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000111111111111111111011111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111111111111111111111110011111111111111111100000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111100111111111111111111100000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101101111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111001111111111111111111000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000111111111111111111111111111111111111111111110111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111111111111111111111111110011111111111111111110000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000001111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111000011111111111111111111111111111111100111111111111111111110000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000001111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111110111111111111111111111111111111111111111111111111111111111111111111111111111000111110000000110011111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111111111000111111111111111111111111111111111111111110000111111111111111111111111111111111000111111111111111111100000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000011111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111110111111111111111111111111111111111000111111111111111111111111111111111111100011111111111111111001111111111111111111111111111111111111111111111111111111110000001111111111111111111111111111111111111100000001111111111111111111111111111111111111000011111111111111111111111111111111110011111111111111111111000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000011111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111110111111111111111111111111111111100000011111111111111111111111111111111110000111111111111111111101111111111111111111111111111111111111111111111111111111000011100111111111111111111111111111111111100001111100111111111111111111111111111111111100001111111111111111111111111111111111100111111111111111111111000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000111111111111111110111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111011111111111111111111111111100000110011111111111111111111111111111111000001111111111111111111100111111111111111111111111111111111111111111111111111000001111110011111111111111111111111111111110000011111100011111111111111111111111111111110000111111111111111111111111111111111111001111111111111111111110000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111001111111111111111111111110000011111100111111111111111111111111111100001111111111111111111111110011111111111111111111111111111111111111111111111110000111111111000111111111111111111111111111000001111111110001111111111111111111111111110000011111111111111111111111111111111111100011111111111111111111100000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111111111111000011111111100011111111111111111111111110000111111111111111111111111111001111111111111111111111100011111111111111111110000111111111111100001111111111111111111111000001111111111111100011111111111111111111111000001111111111111111111111111111111111111000111111111111111111111100000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000001111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000111111111111100000001111111111111000111111111111111111100000001111111111111111111111111111100001111111111111111110000001111111111110000000101111111111111111000011111111111111111000000011111111111111110000111111111111111110000000111111111111111111111111111111111111111001111111111111111111111000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000001111111111111111000011111011111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000001111111111111111110000011111111110000000011111111111111111111111111111111111000000011111111000000111100000100000000000011111111111111111111110000000000000000000000111111111111111111111100000000111110000000001111111111111111111111111111111111111111100011111111111111111111110000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000001111111111111111000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000011111111111111111111111100000000000000000011111111111111111111111111111111111111111000000000000000011111111000000000000111111111111111111111111111110000000000000001111111111111111111111111111100000000000000011111111111111111111111111111111111111111111000111111111111111111111110000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000001111111111111111100111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000001111111111111111111111111111100000000001111111111111111111111111111111111111111111111111100000000011111111111110011111111111111111111111111111111111111111100001111111111111111111111111111111111111111111000111111111111111111111111111111111111111111111100001111111111111111111111000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000001111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111111111111110000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111111111111111110000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111111111111111100000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111111111111111111000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111111111111100000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111111111111111111100000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111111111111111110000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111111111111111111100000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111111111111111111000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000001111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000011111111111000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111110000000001111111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000111111111111111111111111111111111111111111111111111111111000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111100011111011111111100011100011111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000001111111111111111110111111111111111111111111111111100000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011011111111111000111111111111111000111111111111111000111111111110000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000011111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000001111111111111111111111111111111111111111111100000000000001111111111111111111111111111000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111100000001111111111000111111111111111001111111111111111000111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000011111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000001111111111111111111111111111111111111111100000000111111111111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111111111111111111100000011111100011111111111111111100100001111111111000111111111111111000111111111111111000111111111000011110000011111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000011111111111111111111111111111111111111000000001111111111111111111111111111111111111111111111111111111111111111000000000000000000011111111111111111111111111111111111111111111100000000011111100011111111111111111000111000111111111000011111111111111100011111111111111000111111110001111111110111111110000000011111111111111111111111111111111111111111111111111111111111111111111111111111110000000111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000111111111111111111111111111111111111000000111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000111111111111111111111111111111111111111000011100011111100011111111111111111000111000111111111100001111111111111100011111111111111000111111110001111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000111111111111111111111111111111111100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000011111111111111111111111111111110001111111111111100011111111111111110001111100011111111110000011111111111100000111111111111000111111100011111111111111111100011110000111111111111111111111111111111111111111111111111111111111111111111111100000001111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000001111111111111111111111111111111100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000111111111111111111111100011111111111111100011111111111111110011111100011111111111000000111111111111000000111111111000111111100011111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000001111111111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000111111111111111111000111111111111111100011111111111111110011111110011111111111111000001111111111111000011111111000111111100011111111111111111100011111111111111111111111111111111111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000001111111111111111111111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111111100011111111111111100011111111001111111111111110000111111111111100001111111000111111100011111111111111111100011111111111111111111111111111111111111111111111111111111111110000000000011111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000001111111111111111111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111111111100011111111111111100011111110001111111111111111010111111111111110001111111000111111100011111111111111111110001111111111111111111111111111111111111111111111111111110000000000011111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000001111111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111111111100011111111111111100011111100001111111111111111000111111111111111001111111000111111100011111111111111111111000111111111111111111111111111111111111111111111110000000000111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000011111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111100011111111111111000000000000001111111111111111000111111111111111000111111000111111100011111111111111111111110011111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000011111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111100011111111111111000000000000000111111111111111000111111111111111000111111000111111100011111111111111111111111000111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000011111111111111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111100011111111111110000111111111000111111111111110001111111101111110001111111000111111110001111111111111111111111100011111111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000011111111111111011110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111111111100011111111111110001111111111100011111000000000011111111000000000001111111000111111110000111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000011111111111111000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100001111111111111111100011111111111110011111111111110011111100000000111111111000000000011111111000111111111000011111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000011111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111111111100001100001111110011111111111111111111111111111111111111111000011111111111100111111111100001111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000001111111111111111001111111111111111111111111111111111111100000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111110001111111111111111100000000001111110111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000001111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111000111111100011111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000111111100111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000001111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111100011110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000001111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000001111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000011111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000011111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000011111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000011111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000011111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000001111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111110011111100000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000")
);

signal bCoord_X : integer := 0;-- offset from start position 
signal bCoord_Y : integer := 0;

signal drawing_X : std_logic := '0';
signal drawing_Y : std_logic := '0';
	
signal objectEndX : integer;
signal objectEndY : integer;

begin

-- Calculate object end boundaries
objectEndX	<= object_X_size+ObjectStartX;
objectEndY	<= object_Y_size+ObjectStartY;

-- Signals drawing_X[Y] are active when obects coordinates are being crossed

-- test if ooCoord is in the rectangle defined by Start and End 
	drawing_X	<= '1' when  (oCoord_X  >= ObjectStartX) and  (oCoord_X < objectEndX) else '0';
    drawing_Y	<= '1' when  (oCoord_Y  >= ObjectStartY) and  (oCoord_Y < objectEndY) else '0';

-- calculate offset from start corner 
	bCoord_X 	<= (oCoord_X - ObjectStartX) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 
	bCoord_Y 	<= (oCoord_Y - ObjectStartY) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 


process ( RESETn, CLK)

  		
   begin
	if RESETn = '0' then
	    mVGA_RGB	<=  (others => '0') ; 	
		drawing_request	<=  '0' ;

		elsif rising_edge(CLK) then
			mVGA_RGB	<=  object_colors(bCoord_Y , bCoord_X);	--get from colors table 
			drawing_request	<= object(bCoord_Y , bCoord_X) and drawing_X and drawing_Y ; -- get from mask table if inside rectangle  
	end if;

  end process;

		
end behav;
