library IEEE;
use IEEE.STD_LOGIC_1164.all;



entity middle_layer_draw is
port 	(
		--////////////////////	Clock Input	 	////////////////////	
	   CLK  					: in std_logic;
		RESETn				: in std_logic;
		oCoord_X				: in integer;
		oCoord_Y				: in integer;
		random				: in std_logic_vector(1 downto 0);
		endOfFrame			: in std_logic;
		space_was_pressed : in std_logic ;
		game_over			: in std_logic ;
		drawing_request	: out std_logic ;
		mVGA_RGB 			: out std_logic_vector(7 downto 0) 
	);
end entity;

architecture behave of middle_layer_draw is 


	signal sigSpaceWasPressed : std_logic := '0';
	signal sigGameOver : std_logic := '0';
	signal sig_draw_req : std_logic := '0';
	signal sig_draw_data: std_logic_vector (7 downto 0);
	
	constant Draw_Size_X : integer := 200;
	constant Draw_Size_Y : integer := 150;
	
	type ram_array is array(0 to Draw_Size_Y - 1 , 0 to Draw_Size_X - 1) of std_logic_vector(7 downto 0);
	type mask_array is array(0 to Draw_Size_Y - 1, 0 to Draw_Size_X - 1) of std_logic;
	
	signal bCoord_X : integer := 0;-- offset from start position 
	signal bCoord_Y : integer := 0;

	signal drawing_X : std_logic := '0';
	signal drawing_Y : std_logic := '0';
	
	constant ObjectStartX : integer := 214;
	constant objectStartY : integer := 160;

	--		
	signal objectEndX : integer;
	signal objectEndY : integer;
	
	signal sig_color : ram_array;
	signal sig_mask : mask_array;
	
	constant logo1_Colors : ram_array := (
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"92",x"92",x"b6",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"92",x"6d",x"92",x"b6",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"6d",x"6d",x"24",x"6d",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"92",x"92",x"92",x"b6",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"92",x"6d",x"24",x"00",x"49",x"6d",x"92",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"6d",x"6d",x"6d",x"92",x"b6",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"b6",x"92",x"6d",x"49",x"24",x"49",x"24",x"6d",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"b6",x"92",x"6d",x"49",x"25",x"49",x"6d",x"92",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"92",x"49",x"24",x"24",x"b6",x"00",x"49",x"6d",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"49",x"00",x"00",x"24",x"49",x"6d",x"92",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"6d",x"49",x"00",x"6d",x"ff",x"24",x"24",x"6d",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"6d",x"24",x"00",x"00",x"00",x"24",x"6d",x"6d",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"b6",x"92",x"92",x"92",x"92",x"6d",x"6d",x"49",x"24",x"00",x"b6",x"ff",x"49",x"00",x"49",x"92",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"6d",x"24",x"00",x"25",x"00",x"00",x"48",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"da",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"49",x"24",x"00",x"24",x"ff",x"ff",x"6d",x"00",x"49",x"6d",x"92",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"6d",x"24",x"25",x"97",x"00",x"00",x"24",x"49",x"49",x"6d",x"6d",x"71",x"91",x"91",x"92",x"92",x"71",x"71",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b7",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"92",x"92",x"92",x"92",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b7",x"db",x"db",x"db",x"ff",x"db",x"b6",x"92",x"6d",x"6d",x"69",x"49",x"49",x"49",x"24",x"24",x"00",x"92",x"ff",x"ff",x"b6",x"00",x"24",x"6d",x"92",x"92",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b7",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"24",x"25",x"ff",x"25",x"00",x"00",x"24",x"45",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"b6",x"6d",x"6d",x"6d",x"6d",x"92",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"b6",x"db",x"db",x"db",x"db",x"b6",x"6d",x"49",x"29",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"bb",x"ff",x"ff",x"db",x"00",x"24",x"49",x"6d",x"92",x"92",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"b6",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"b2",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"49",x"00",x"49",x"ff",x"b2",x"00",x"00",x"04",x"24",x"24",x"45",x"45",x"45",x"45",x"49",x"48",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6e",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"92",x"6d",x"49",x"24",x"49",x"6d",x"92",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"b6",x"db",x"db",x"b6",x"92",x"6d",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"ff",x"ff",x"ff",x"ff",x"24",x"00",x"24",x"49",x"6d",x"6d",x"92",x"b6",x"b6",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"91",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"49",x"00",x"45",x"ff",x"fa",x"8e",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"04",x"00",x"04",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"92",x"6d",x"49",x"00",x"00",x"20",x"49",x"6d",x"92",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"b6",x"b6",x"b6",x"92",x"6d",x"49",x"00",x"20",x"69",x"00",x"00",x"00",x"00",x"00",x"92",x"ff",x"ff",x"ff",x"ff",x"49",x"00",x"24",x"24",x"49",x"6d",x"6d",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"49",x"00",x"25",x"fb",x"d6",x"d6",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"92",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"92",x"6d",x"49",x"24",x"24",x"92",x"00",x"24",x"49",x"6d",x"92",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b7",x"92",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"92",x"b6",x"b6",x"92",x"6d",x"24",x"00",x"60",x"f6",x"df",x"ff",x"fb",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"6d",x"00",x"00",x"00",x"24",x"49",x"49",x"6d",x"92",x"b6",x"b6",x"b6",x"92",x"6d",x"6d",x"49",x"24",x"48",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"28",x"49",x"6d",x"92",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"00",x"00",x"fb",x"d5",x"f6",x"fb",x"6e",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"49",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"6d",x"92",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"6d",x"49",x"49",x"00",x"49",x"db",x"00",x"00",x"45",x"49",x"6d",x"92",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"91",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"6d",x"92",x"92",x"6d",x"49",x"04",x"20",x"80",x"ee",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"24",x"00",x"00",x"00",x"00",x"49",x"6d",x"6d",x"92",x"92",x"92",x"6d",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"49",x"6d",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"24",x"00",x"b7",x"fa",x"d1",x"f6",x"fb",x"d6",x"92",x"6d",x"8d",x"92",x"b2",x"d6",x"db",x"db",x"fb",x"fb",x"db",x"db",x"92",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"6d",x"92",x"b6",x"db",x"db",x"db",x"db",x"b6",x"92",x"6d",x"49",x"49",x"24",x"00",x"92",x"ff",x"29",x"00",x"24",x"49",x"49",x"6d",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"6d",x"92",x"92",x"6d",x"49",x"00",x"20",x"c4",x"c4",x"f6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"92",x"49",x"00",x"00",x"24",x"6d",x"6d",x"6d",x"6d",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"49",x"6d",x"92",x"b6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"6d",x"24",x"00",x"6e",x"ff",x"d0",x"d0",x"f5",x"fa",x"fb",x"fb",x"fb",x"fb",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"ff",x"ff",x"d7",x"49",x"00",x"00",x"00",x"00",x"49",x"96",x"b7",x"db",x"db",x"db",x"b7",x"92",x"25",x"00",x"00",x"00",x"24",x"6d",x"92",x"b6",x"db",x"db",x"db",x"db",x"b6",x"92",x"6d",x"49",x"24",x"00",x"00",x"db",x"ff",x"72",x"00",x"00",x"24",x"49",x"6d",x"92",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"24",x"00",x"69",x"92",x"b6",x"b6",x"96",x"b2",x"b2",x"b2",x"b2",x"b6",x"8e",x"00",x"24",x"6d",x"6d",x"6d",x"49",x"24",x"00",x"40",x"e4",x"e0",x"c9",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"6d",x"04",x"49",x"6d",x"6d",x"49",x"24",x"24",x"00",x"00",x"00",x"6e",x"b6",x"b7",x"b7",x"b6",x"92",x"25",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"49",x"92",x"b7",x"b7",x"b6",x"92",x"49",x"00",x"00",x"00",x"24",x"49",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"6d",x"24",x"00",x"24",x"fb",x"d5",x"ac",x"f0",x"f0",x"f5",x"f5",x"f5",x"f5",x"f5",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f5",x"fa",x"da",x"6e",x"00",x"49",x"b2",x"db",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"fa",x"d6",x"92",x"00",x"00",x"00",x"48",x"6d",x"92",x"b6",x"db",x"db",x"b6",x"92",x"6d",x"49",x"00",x"00",x"00",x"24",x"ff",x"ff",x"bb",x"00",x"00",x"00",x"00",x"24",x"6d",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"71",x"49",x"00",x"00",x"db",x"ff",x"fe",x"fa",x"fa",x"fa",x"fa",x"fa",x"d6",x"ff",x"db",x"00",x"00",x"49",x"6d",x"6d",x"49",x"24",x"00",x"80",x"e0",x"e0",x"e0",x"f2",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"b6",x"00",x"48",x"48",x"49",x"24",x"00",x"00",x"00",x"69",x"b6",x"fb",x"fa",x"fa",x"f6",x"fa",x"fa",x"d7",x"6e",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"92",x"db",x"fe",x"fa",x"fa",x"f6",x"fb",x"db",x"92",x"25",x"00",x"00",x"49",x"6d",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"49",x"00",x"00",x"b6",x"ff",x"b1",x"ac",x"f0",x"f0",x"f0",x"f0",x"f0",x"f0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"fa",x"fb",x"92",x"d7",x"fa",x"f5",x"f1",x"ec",x"f0",x"f0",x"f0",x"f5",x"f5",x"fa",x"fb",x"b2",x"20",x"00",x"24",x"49",x"6e",x"92",x"b6",x"b6",x"92",x"6d",x"49",x"24",x"49",x"6d",x"6d",x"b6",x"ff",x"ff",x"df",x"92",x"6d",x"49",x"00",x"20",x"49",x"6d",x"96",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"6d",x"45",x"00",x"25",x"ff",x"f9",x"f9",x"f9",x"f5",x"f5",x"f4",x"f0",x"ad",x"db",x"b7",x"00",x"24",x"49",x"6d",x"49",x"49",x"00",x"20",x"c4",x"e0",x"e0",x"e0",x"e5",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"8d",x"00",x"24",x"28",x"25",x"00",x"00",x"00",x"6d",x"fb",x"fe",x"f9",x"f5",x"f0",x"f0",x"f0",x"f5",x"f6",x"fb",x"92",x"00",x"00",x"00",x"00",x"49",x"d7",x"ff",x"fa",x"f9",x"f4",x"f0",x"f0",x"f1",x"fa",x"fb",x"b6",x"24",x"00",x"24",x"6d",x"92",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"92",x"49",x"24",x"00",x"29",x"ff",x"fa",x"ad",x"ac",x"cc",x"f0",x"f0",x"f0",x"f0",x"f0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f6",x"fb",x"f6",x"ed",x"e8",x"e8",x"ec",x"ec",x"f0",x"f0",x"f4",x"f4",x"f4",x"f5",x"fa",x"92",x"00",x"00",x"24",x"6d",x"6d",x"92",x"92",x"6d",x"6d",x"24",x"24",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"d6",x"69",x"00",x"24",x"49",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"24",x"00",x"6e",x"fe",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"ec",x"88",x"db",x"6e",x"00",x"24",x"49",x"6d",x"49",x"24",x"00",x"40",x"c4",x"e0",x"e4",x"e0",x"e0",x"f2",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ae",x"20",x"00",x"24",x"24",x"24",x"00",x"00",x"6e",x"fb",x"fe",x"f9",x"f4",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"f6",x"fb",x"49",x"00",x"00",x"45",x"db",x"fe",x"f9",x"f4",x"f4",x"f0",x"ec",x"ec",x"ec",x"ec",x"f1",x"fb",x"92",x"00",x"00",x"49",x"92",x"b6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"92",x"49",x"24",x"00",x"00",x"72",x"ff",x"da",x"8d",x"88",x"a8",x"cc",x"cc",x"f0",x"f0",x"f0",x"f0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"ec",x"f1",x"ec",x"e8",x"e8",x"e8",x"ec",x"f0",x"f0",x"f4",x"f4",x"f4",x"f0",x"f0",x"f5",x"fb",x"49",x"00",x"24",x"49",x"6d",x"6d",x"6d",x"6d",x"49",x"24",x"00",x"92",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"f6",x"a5",x"20",x"04",x"49",x"6d",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"49",x"00",x"00",x"b6",x"f9",x"f4",x"f4",x"f4",x"f4",x"f0",x"ec",x"ec",x"ad",x"ff",x"49",x"00",x"24",x"49",x"49",x"49",x"04",x"00",x"60",x"e4",x"e0",x"e4",x"e0",x"e0",x"c5",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"d2",x"60",x"00",x"04",x"24",x"24",x"00",x"00",x"49",x"fb",x"fe",x"f8",x"f4",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"f6",x"b6",x"00",x"04",x"b7",x"ff",x"f8",x"f4",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"f1",x"db",x"25",x"00",x"49",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"92",x"6d",x"49",x"24",x"00",x"00",x"96",x"ff",x"fb",x"b1",x"8d",x"88",x"88",x"ac",x"d0",x"f0",x"f0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"ec",x"f0",x"f0",x"f4",x"f4",x"f4",x"f4",x"f0",x"ec",x"f6",x"b2",x"00",x"00",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"00",x"24",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"f6",x"e5",x"c0",x"40",x"00",x"24",x"6d",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"49",x"00",x"00",x"db",x"f9",x"f4",x"f4",x"f4",x"f4",x"f0",x"ec",x"c8",x"b1",x"db",x"00",x"00",x"24",x"49",x"49",x"49",x"00",x"00",x"a0",x"e0",x"e0",x"e4",x"e0",x"e0",x"c0",x"f6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"f2",x"84",x"20",x"00",x"04",x"00",x"20",x"00",x"00",x"b6",x"fe",x"f8",x"f8",x"f4",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"cd",x"db",x"25",x"6e",x"ff",x"f9",x"f8",x"f4",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"cc",x"fa",x"6e",x"00",x"24",x"6d",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"6d",x"49",x"24",x"00",x"00",x"04",x"96",x"ff",x"ff",x"ff",x"d6",x"b2",x"8d",x"ac",x"d0",x"f0",x"f0",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"ec",x"e8",x"e8",x"a4",x"a4",x"a8",x"cc",x"f0",x"f0",x"f4",x"f4",x"f4",x"f4",x"f0",x"ec",x"d1",x"db",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"49",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ed",x"e0",x"e0",x"80",x"00",x"24",x"49",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"db",x"b6",x"6d",x"49",x"00",x"25",x"ff",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"ec",x"88",x"d6",x"b7",x"00",x"00",x"24",x"49",x"49",x"24",x"00",x"20",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"a5",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"f6",x"a5",x"60",x"00",x"00",x"00",x"00",x"00",x"00",x"6e",x"ff",x"f8",x"f8",x"f4",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"c8",x"da",x"92",x"db",x"f9",x"f8",x"f8",x"f4",x"f0",x"ec",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"c8",x"d6",x"96",x"00",x"24",x"6d",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"44",x"24",x"00",x"00",x"00",x"6e",x"db",x"ff",x"ff",x"ff",x"fb",x"d6",x"d0",x"f0",x"f0",x"f4",x"f4",x"f4",x"f4",x"f0",x"ec",x"ec",x"e8",x"84",x"64",x"69",x"8d",x"cc",x"ec",x"f0",x"f4",x"f4",x"f4",x"f4",x"ec",x"ec",x"cc",x"fb",x"25",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"db",x"ff",x"ff",x"ff",x"ff",x"f6",x"c0",x"e0",x"e0",x"c0",x"40",x"00",x"24",x"6d",x"92",x"db",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"24",x"00",x"6d",x"fe",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"ec",x"88",x"db",x"6e",x"00",x"24",x"24",x"49",x"49",x"24",x"00",x"60",x"e4",x"e0",x"e0",x"e0",x"e0",x"c0",x"ad",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"cd",x"80",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"db",x"f9",x"f4",x"f4",x"f4",x"f0",x"ec",x"ec",x"c8",x"c4",x"e8",x"ec",x"ec",x"e8",x"c8",x"d6",x"ff",x"fa",x"f8",x"f8",x"f4",x"f4",x"f0",x"ec",x"c8",x"c4",x"e8",x"ec",x"ec",x"ec",x"c8",x"b1",x"bb",x"00",x"24",x"6d",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"24",x"24",x"00",x"00",x"00",x"25",x"92",x"b7",x"db",x"ff",x"ff",x"da",x"f0",x"f0",x"f0",x"f4",x"f4",x"f4",x"f0",x"ec",x"ec",x"c8",x"64",x"b6",x"ff",x"fb",x"d6",x"f0",x"f0",x"f4",x"f4",x"f4",x"f0",x"f0",x"ec",x"c8",x"fb",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"db",x"ff",x"ff",x"ff",x"ff",x"d6",x"c5",x"e0",x"e0",x"e0",x"60",x"00",x"24",x"6d",x"92",x"b6",x"db",x"ff",x"db",x"b6",x"92",x"49",x"24",x"00",x"b6",x"fa",x"f4",x"f4",x"f4",x"f4",x"f0",x"ec",x"c8",x"8d",x"ff",x"29",x"00",x"24",x"49",x"49",x"28",x"20",x"00",x"84",x"e0",x"e0",x"e0",x"e0",x"e0",x"c5",x"b6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ad",x"40",x"00",x"00",x"00",x"20",x"00",x"00",x"69",x"ff",x"f8",x"f8",x"f4",x"f4",x"f0",x"ec",x"ec",x"84",x"84",x"e8",x"e8",x"e8",x"ec",x"a8",x"d6",x"ff",x"f9",x"f4",x"f4",x"f4",x"f0",x"ec",x"ec",x"a8",x"84",x"c8",x"ec",x"ec",x"ec",x"c8",x"ad",x"db",x"00",x"24",x"6d",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"6d",x"4d",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"24",x"24",x"04",x"00",x"00",x"00",x"00",x"00",x"25",x"6e",x"db",x"ff",x"f0",x"f0",x"f0",x"f4",x"f4",x"f0",x"f0",x"ec",x"e8",x"84",x"b2",x"ff",x"ff",x"ff",x"ff",x"d1",x"f0",x"f4",x"f4",x"f4",x"f0",x"f0",x"ec",x"a8",x"fb",x"49",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"a9",x"e0",x"e4",x"e0",x"a0",x"00",x"20",x"49",x"92",x"b6",x"db",x"db",x"db",x"b6",x"92",x"49",x"00",x"00",x"db",x"f5",x"f4",x"f4",x"f4",x"f4",x"f0",x"ec",x"c8",x"b1",x"db",x"00",x"00",x"24",x"49",x"49",x"24",x"00",x"00",x"a4",x"e0",x"e4",x"e0",x"e0",x"e4",x"a9",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"8d",x"00",x"00",x"20",x"20",x"00",x"00",x"00",x"b7",x"fa",x"f4",x"f8",x"f4",x"f0",x"f0",x"e8",x"c8",x"89",x"d7",x"f1",x"e8",x"e8",x"e8",x"a4",x"da",x"fa",x"f8",x"f8",x"f4",x"f0",x"f0",x"ec",x"e8",x"88",x"d6",x"f1",x"ec",x"ec",x"ec",x"a4",x"d6",x"b6",x"00",x"24",x"6d",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"4d",x"28",x"00",x"24",x"24",x"44",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"db",x"f9",x"f0",x"f0",x"f4",x"f4",x"f0",x"f0",x"ec",x"c8",x"69",x"ff",x"db",x"6e",x"6e",x"fb",x"f5",x"f0",x"f0",x"f4",x"f0",x"f0",x"ec",x"ec",x"88",x"ff",x"49",x"00",x"00",x"6d",x"d7",x"db",x"db",x"92",x"25",x"00",x"00",x"49",x"ff",x"ff",x"df",x"ff",x"ff",x"df",x"92",x"c4",x"e0",x"e4",x"c4",x"20",x"00",x"29",x"6d",x"b6",x"ba",x"db",x"db",x"92",x"6d",x"24",x"00",x"28",x"fb",x"f0",x"f4",x"f4",x"f4",x"f0",x"f0",x"ec",x"84",x"d6",x"b6",x"00",x"00",x"24",x"49",x"49",x"24",x"00",x"40",x"e4",x"e4",x"e0",x"e0",x"e0",x"c4",x"92",x"bf",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"6e",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"ff",x"f8",x"f4",x"f4",x"f4",x"f0",x"ec",x"ec",x"a4",x"b2",x"ff",x"f1",x"e4",x"e8",x"c8",x"a8",x"ff",x"f9",x"f4",x"f4",x"f4",x"f0",x"ec",x"ec",x"c8",x"8d",x"ff",x"f6",x"e8",x"ec",x"e8",x"88",x"db",x"92",x"00",x"24",x"6d",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"6d",x"49",x"00",x"00",x"00",x"00",x"24",x"24",x"25",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"b6",x"f5",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"a4",x"d6",x"ff",x"49",x"00",x"00",x"d7",x"f5",x"f0",x"f0",x"f4",x"f0",x"f0",x"ec",x"e8",x"ad",x"ff",x"05",x"25",x"b6",x"ff",x"fe",x"fe",x"fa",x"fb",x"d7",x"25",x"00",x"6d",x"ff",x"9f",x"9b",x"b6",x"ff",x"df",x"9b",x"a9",x"e0",x"e0",x"e0",x"60",x"00",x"24",x"6d",x"92",x"b6",x"db",x"b6",x"92",x"6d",x"24",x"00",x"6d",x"fa",x"f0",x"f4",x"f4",x"f4",x"f0",x"ec",x"ec",x"84",x"fb",x"6e",x"00",x"00",x"24",x"49",x"49",x"24",x"00",x"60",x"e4",x"e0",x"e0",x"e0",x"e0",x"c9",x"97",x"bf",x"ff",x"ff",x"ff",x"fb",x"db",x"ff",x"ff",x"ff",x"ff",x"8d",x"00",x"00",x"00",x"00",x"00",x"00",x"69",x"fb",x"f4",x"f4",x"f4",x"f4",x"f0",x"ec",x"e8",x"a4",x"db",x"ff",x"ec",x"e8",x"e8",x"c8",x"ad",x"ff",x"f5",x"f4",x"f4",x"f0",x"f0",x"ec",x"e8",x"a4",x"b2",x"ff",x"f1",x"e8",x"e8",x"e8",x"a8",x"df",x"6d",x"00",x"24",x"6d",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"6d",x"49",x"00",x"24",x"96",x"00",x"00",x"00",x"00",x"24",x"24",x"28",x"49",x"49",x"44",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"d7",x"f5",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"ec",x"84",x"fb",x"92",x"00",x"00",x"00",x"db",x"f5",x"f0",x"f4",x"f0",x"f0",x"ec",x"ec",x"c8",x"b1",x"db",x"25",x"d7",x"fe",x"f9",x"f4",x"f4",x"f4",x"f5",x"fa",x"92",x"00",x"92",x"bf",x"5b",x"5b",x"72",x"d2",x"ff",x"7b",x"92",x"c0",x"e0",x"e0",x"a0",x"00",x"00",x"49",x"92",x"b6",x"b6",x"b6",x"92",x"49",x"00",x"00",x"b6",x"fa",x"f0",x"f4",x"f4",x"f0",x"f0",x"ec",x"c8",x"a9",x"ff",x"25",x"00",x"24",x"24",x"49",x"24",x"00",x"00",x"a0",x"e0",x"e0",x"e0",x"e0",x"c0",x"ae",x"7b",x"df",x"ff",x"ff",x"fb",x"b2",x"76",x"df",x"ff",x"ff",x"ff",x"92",x"00",x"00",x"00",x"24",x"00",x"00",x"b6",x"fa",x"f4",x"f4",x"f4",x"f0",x"ec",x"e8",x"e8",x"88",x"ff",x"fa",x"e8",x"e8",x"e8",x"a4",x"b6",x"fe",x"f4",x"f4",x"f4",x"f0",x"f0",x"ec",x"e8",x"84",x"db",x"ff",x"cd",x"e8",x"e8",x"c8",x"ad",x"ff",x"25",x"00",x"49",x"6d",x"b6",x"db",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"92",x"6d",x"45",x"00",x"b6",x"bf",x"7b",x"2d",x"00",x"00",x"00",x"04",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"25",x"fb",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"c8",x"88",x"db",x"25",x"00",x"00",x"29",x"ff",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"a8",x"d6",x"b7",x"d7",x"ff",x"f9",x"f8",x"f4",x"f4",x"f0",x"ec",x"d1",x"db",x"00",x"76",x"7b",x"5b",x"5f",x"7b",x"89",x"d2",x"7b",x"77",x"c5",x"e0",x"e0",x"c4",x"40",x"00",x"29",x"6d",x"92",x"b6",x"92",x"6d",x"24",x"00",x"00",x"db",x"f5",x"f4",x"f4",x"f0",x"f0",x"ec",x"ec",x"c8",x"b2",x"db",x"00",x"00",x"24",x"24",x"49",x"24",x"00",x"20",x"c4",x"e0",x"e0",x"e4",x"e0",x"c4",x"92",x"7f",x"ff",x"ff",x"f6",x"a5",x"8d",x"7b",x"7b",x"bf",x"ff",x"ff",x"b6",x"00",x"00",x"00",x"00",x"00",x"00",x"db",x"f9",x"f4",x"f4",x"f4",x"f0",x"ec",x"e8",x"c4",x"ad",x"ff",x"f6",x"e4",x"e8",x"e4",x"a4",x"da",x"fa",x"f0",x"f0",x"f0",x"f0",x"ec",x"e8",x"e8",x"88",x"ff",x"fb",x"c8",x"e8",x"e8",x"a4",x"b2",x"db",x"00",x"00",x"49",x"92",x"b6",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"6d",x"49",x"24",x"04",x"db",x"9b",x"5b",x"5b",x"2e",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"6d",x"fb",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"e8",x"a4",x"b1",x"db",x"24",x"00",x"00",x"6e",x"fa",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"e8",x"88",x"db",x"db",x"fa",x"f5",x"f4",x"f4",x"f4",x"f0",x"ec",x"ec",x"ac",x"fb",x"49",x"2e",x"7b",x"5b",x"3f",x"5f",x"92",x"a4",x"92",x"7b",x"ae",x"e0",x"e0",x"c4",x"80",x"00",x"24",x"4d",x"92",x"92",x"92",x"6d",x"24",x"00",x"49",x"fb",x"f4",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"a8",x"d6",x"97",x"00",x"00",x"24",x"49",x"49",x"24",x"00",x"60",x"e4",x"e0",x"e0",x"e0",x"e0",x"a9",x"7b",x"9f",x"ff",x"ed",x"c4",x"a5",x"76",x"5f",x"5b",x"7b",x"df",x"ff",x"db",x"00",x"00",x"00",x"00",x"00",x"25",x"ff",x"f4",x"f4",x"f0",x"f0",x"f0",x"ec",x"e8",x"a4",x"d6",x"ff",x"ed",x"e4",x"e8",x"e4",x"84",x"ff",x"f5",x"f0",x"f0",x"f0",x"ec",x"ec",x"e8",x"c8",x"ad",x"ff",x"f6",x"e8",x"e8",x"e8",x"84",x"da",x"96",x"00",x"00",x"49",x"92",x"b6",x"db",x"db",x"db",x"b6",x"b6",x"92",x"92",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"24",x"00",x"49",x"ff",x"bf",x"5b",x"5b",x"7f",x"77",x"29",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"b2",x"fa",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"e8",x"84",x"d6",x"b7",x"00",x"00",x"00",x"b6",x"f6",x"f0",x"f0",x"f0",x"f0",x"ec",x"e8",x"c8",x"8d",x"ff",x"ff",x"f5",x"f4",x"f4",x"f0",x"f0",x"f0",x"ec",x"ec",x"a8",x"da",x"4a",x"00",x"77",x"5f",x"3f",x"5b",x"97",x"a9",x"89",x"9b",x"76",x"c5",x"e0",x"e4",x"80",x"20",x"04",x"49",x"8e",x"92",x"6d",x"49",x"00",x"00",x"8e",x"fa",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"e8",x"88",x"fb",x"6e",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"80",x"e0",x"e0",x"e0",x"e0",x"c4",x"92",x"7f",x"bb",x"c9",x"c0",x"c0",x"ae",x"7f",x"3b",x"3b",x"5f",x"9f",x"df",x"db",x"00",x"00",x"00",x"00",x"00",x"6d",x"fa",x"f4",x"f4",x"f0",x"f0",x"ec",x"e8",x"e8",x"84",x"db",x"fb",x"e8",x"e4",x"e8",x"c4",x"8d",x"ff",x"f4",x"f0",x"f0",x"f0",x"ec",x"e8",x"e8",x"a4",x"d2",x"ff",x"f1",x"e8",x"e8",x"e8",x"88",x"ff",x"6e",x"00",x"24",x"49",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"6d",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"b6",x"92",x"6d",x"6d",x"49",x"24",x"00",x"92",x"ff",x"bf",x"5b",x"5b",x"5b",x"5f",x"7b",x"2d",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"db",x"f5",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"e8",x"88",x"ff",x"6e",x"00",x"00",x"00",x"db",x"f5",x"f0",x"f0",x"f0",x"ec",x"ec",x"e8",x"a8",x"b2",x"ff",x"ff",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"e8",x"88",x"da",x"6e",x"00",x"29",x"5b",x"3b",x"5b",x"5b",x"92",x"a5",x"92",x"7b",x"89",x"e0",x"e0",x"a0",x"20",x"00",x"49",x"6d",x"6d",x"6d",x"49",x"00",x"00",x"b6",x"f9",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"c8",x"8d",x"ff",x"25",x"00",x"24",x"49",x"49",x"24",x"00",x"20",x"80",x"c0",x"c0",x"c0",x"e0",x"a9",x"77",x"7b",x"a9",x"c0",x"e0",x"c9",x"97",x"5b",x"5b",x"5f",x"5b",x"5b",x"9f",x"df",x"24",x"00",x"00",x"00",x"00",x"b6",x"f9",x"f4",x"f0",x"f0",x"f0",x"ec",x"e8",x"c4",x"89",x"ff",x"f6",x"e4",x"e4",x"e8",x"a4",x"b6",x"fa",x"f0",x"f0",x"f0",x"ec",x"ec",x"e8",x"e8",x"84",x"db",x"ff",x"ec",x"e8",x"e8",x"c4",x"8d",x"ff",x"25",x"00",x"24",x"49",x"92",x"92",x"b6",x"92",x"92",x"92",x"6d",x"49",x"49",x"49",x"49",x"6d",x"92",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"b6",x"92",x"6d",x"6d",x"49",x"24",x"00",x"24",x"db",x"ff",x"df",x"7b",x"5b",x"3b",x"3b",x"5b",x"7b",x"52",x"04",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"fb",x"f1",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"e8",x"89",x"ff",x"45",x"00",x"00",x"45",x"fb",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"a4",x"d6",x"ff",x"fa",x"f0",x"f0",x"ec",x"f0",x"ec",x"ec",x"e8",x"c8",x"85",x"ff",x"49",x"00",x"00",x"52",x"5f",x"3b",x"5b",x"77",x"a5",x"8d",x"7b",x"92",x"c0",x"e0",x"c0",x"40",x"00",x"24",x"49",x"6d",x"49",x"45",x"00",x"00",x"fb",x"f5",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"c8",x"b1",x"db",x"00",x"00",x"24",x"49",x"49",x"24",x"00",x"20",x"a0",x"c0",x"c0",x"c0",x"e0",x"ad",x"7b",x"72",x"c0",x"e0",x"c0",x"ae",x"5b",x"5b",x"7b",x"5b",x"5b",x"5b",x"7b",x"df",x"49",x"00",x"00",x"00",x"00",x"db",x"f9",x"f0",x"f4",x"f0",x"ec",x"ec",x"e8",x"a4",x"8d",x"ff",x"f1",x"e4",x"e4",x"e4",x"84",x"db",x"fa",x"f0",x"f0",x"f0",x"ec",x"ec",x"e8",x"e8",x"88",x"ff",x"fa",x"c8",x"e8",x"e8",x"a4",x"b2",x"db",x"00",x"00",x"24",x"49",x"6d",x"92",x"92",x"92",x"6d",x"6d",x"49",x"24",x"24",x"00",x"24",x"49",x"49",x"92",x"b6",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"6d",x"6d",x"49",x"24",x"24",x"00",x"49",x"ff",x"ff",x"ff",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"57",x"29",x"00",x"00",x"00",x"04",x"00",x"00",x"00",x"6d",x"fa",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"c8",x"b1",x"db",x"04",x"00",x"00",x"6e",x"fa",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"e8",x"84",x"db",x"ff",x"f5",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"84",x"92",x"df",x"25",x"00",x"00",x"29",x"7b",x"5b",x"5b",x"5b",x"92",x"89",x"92",x"77",x"a5",x"c0",x"c0",x"80",x"00",x"24",x"49",x"49",x"49",x"24",x"00",x"49",x"ff",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"e8",x"a4",x"db",x"b6",x"00",x"00",x"24",x"49",x"49",x"24",x"00",x"40",x"80",x"a0",x"c0",x"e0",x"c0",x"76",x"7b",x"ad",x"e0",x"e0",x"a9",x"97",x"5f",x"5b",x"5b",x"5b",x"5b",x"5b",x"5f",x"9b",x"45",x"00",x"00",x"00",x"45",x"ff",x"f4",x"f0",x"f0",x"f0",x"ec",x"e8",x"e8",x"a4",x"b6",x"ff",x"ed",x"e4",x"e4",x"e4",x"88",x"ff",x"f5",x"f0",x"f0",x"f0",x"ec",x"ec",x"e8",x"c4",x"ad",x"ff",x"f1",x"e4",x"e8",x"e8",x"a4",x"db",x"92",x"00",x"00",x"24",x"49",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"20",x"49",x"6d",x"92",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"db",x"db",x"92",x"6d",x"49",x"49",x"24",x"00",x"00",x"00",x"b6",x"ff",x"ff",x"ff",x"7f",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"57",x"2e",x"00",x"00",x"00",x"00",x"00",x"00",x"92",x"fa",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"e8",x"a4",x"d6",x"b7",x"00",x"00",x"00",x"b6",x"fa",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"c4",x"88",x"ff",x"df",x"f6",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"a4",x"64",x"db",x"96",x"00",x"00",x"00",x"00",x"2e",x"5b",x"3b",x"5b",x"76",x"85",x"89",x"77",x"8d",x"a0",x"c0",x"80",x"20",x"00",x"44",x"49",x"25",x"00",x"00",x"6e",x"fa",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"e8",x"88",x"fb",x"6e",x"00",x"00",x"49",x"49",x"49",x"24",x"00",x"40",x"80",x"a0",x"c0",x"c0",x"a9",x"77",x"77",x"a9",x"e0",x"e0",x"8d",x"7b",x"5b",x"5f",x"5b",x"5b",x"5b",x"5b",x"5f",x"52",x"00",x"00",x"00",x"00",x"8e",x"fe",x"f4",x"f0",x"f0",x"f0",x"ec",x"e8",x"e8",x"a4",x"da",x"ff",x"e8",x"e4",x"e4",x"c4",x"ad",x"ff",x"f5",x"f0",x"f0",x"ec",x"ec",x"e8",x"e8",x"a4",x"d2",x"ff",x"ed",x"e4",x"e8",x"e8",x"84",x"ff",x"6e",x"00",x"00",x"24",x"49",x"69",x"4d",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"4d",x"72",x"00",x"24",x"49",x"6d",x"92",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"49",x"00",x"00",x"00",x"00",x"00",x"49",x"ff",x"ff",x"ff",x"ff",x"bf",x"5f",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5b",x"2e",x"04",x"00",x"00",x"00",x"00",x"db",x"f5",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"e8",x"84",x"fb",x"6e",x"00",x"00",x"00",x"db",x"f5",x"f0",x"f0",x"f0",x"f0",x"ec",x"e8",x"c4",x"b1",x"db",x"b7",x"fa",x"a8",x"e8",x"e8",x"ec",x"c8",x"84",x"64",x"d6",x"ff",x"49",x"00",x"00",x"00",x"00",x"04",x"57",x"5b",x"3b",x"57",x"8e",x"85",x"72",x"52",x"80",x"a0",x"80",x"20",x"00",x"24",x"44",x"24",x"00",x"00",x"b6",x"fa",x"f0",x"f0",x"f0",x"f0",x"ec",x"e8",x"c8",x"89",x"ff",x"49",x"00",x"24",x"49",x"4d",x"49",x"24",x"00",x"40",x"80",x"80",x"a0",x"a0",x"8e",x"5b",x"8d",x"c4",x"e0",x"c5",x"96",x"5b",x"5b",x"5b",x"3b",x"3f",x"5b",x"7b",x"57",x"04",x"00",x"00",x"00",x"00",x"b6",x"fa",x"f0",x"f0",x"f0",x"ec",x"ec",x"e8",x"c4",x"a8",x"ff",x"fa",x"e4",x"e4",x"e4",x"a4",x"d2",x"fa",x"f0",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"84",x"db",x"ff",x"ec",x"e8",x"e8",x"c4",x"ad",x"ff",x"25",x"00",x"00",x"24",x"45",x"49",x"49",x"29",x"24",x"00",x"00",x"00",x"29",x"32",x"7b",x"bf",x"24",x"00",x"24",x"49",x"6d",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"db",x"b6",x"6d",x"49",x"6d",x"6d",x"6d",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"df",x"bf",x"bf",x"bf",x"9f",x"9f",x"97",x"7b",x"5b",x"3b",x"57",x"32",x"25",x"00",x"00",x"25",x"fb",x"f0",x"f0",x"f0",x"f0",x"f0",x"ec",x"e8",x"e8",x"ad",x"df",x"49",x"00",x"00",x"49",x"fb",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"e8",x"a4",x"da",x"b6",x"6e",x"ff",x"ad",x"84",x"80",x"80",x"60",x"68",x"b2",x"ff",x"b7",x"20",x"00",x"00",x"00",x"00",x"00",x"29",x"57",x"3b",x"3b",x"73",x"64",x"69",x"52",x"65",x"80",x"60",x"20",x"00",x"24",x"24",x"24",x"00",x"04",x"fb",x"f5",x"f0",x"f0",x"f0",x"f0",x"ec",x"e8",x"a8",x"b1",x"db",x"00",x"00",x"24",x"49",x"6d",x"49",x"24",x"00",x"20",x"60",x"80",x"80",x"80",x"52",x"56",x"a4",x"e0",x"c0",x"8e",x"7b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5f",x"7b",x"29",x"00",x"00",x"00",x"00",x"00",x"db",x"f5",x"f0",x"f0",x"f0",x"ec",x"ec",x"e8",x"c4",x"ad",x"ff",x"f2",x"e4",x"e4",x"e4",x"84",x"db",x"fa",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e4",x"84",x"ff",x"fa",x"e8",x"e8",x"e8",x"a4",x"b2",x"db",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"4d",x"77",x"7b",x"7b",x"df",x"92",x"00",x"24",x"24",x"49",x"6d",x"b6",x"db",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"db",x"b6",x"6d",x"24",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"ae",x"8e",x"77",x"5b",x"3b",x"37",x"2e",x"04",x"00",x"6d",x"fa",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"e8",x"c4",x"b1",x"db",x"00",x"00",x"00",x"6e",x"fa",x"ec",x"f0",x"f0",x"f0",x"ec",x"ec",x"e8",x"88",x"df",x"6e",x"25",x"db",x"fa",x"b1",x"89",x"89",x"8d",x"d6",x"ff",x"db",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"2e",x"37",x"37",x"57",x"49",x"45",x"2e",x"49",x"60",x"60",x"20",x"00",x"24",x"24",x"20",x"00",x"49",x"fb",x"f0",x"f0",x"f0",x"f0",x"ec",x"e8",x"e8",x"84",x"da",x"b6",x"00",x"00",x"24",x"49",x"6d",x"6d",x"49",x"00",x"20",x"40",x"60",x"60",x"65",x"57",x"6a",x"c0",x"e0",x"a5",x"76",x"5f",x"5b",x"3f",x"5b",x"7b",x"5b",x"5f",x"52",x"00",x"00",x"00",x"00",x"00",x"29",x"ff",x"f4",x"f0",x"f0",x"ec",x"ec",x"e8",x"e8",x"a4",x"b6",x"ff",x"ed",x"e4",x"e4",x"e4",x"88",x"ff",x"f5",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"c4",x"ad",x"ff",x"f1",x"e4",x"e8",x"e4",x"84",x"db",x"92",x"00",x"00",x"00",x"00",x"04",x"24",x"20",x"00",x"00",x"09",x"52",x"7b",x"7b",x"5b",x"7b",x"df",x"db",x"20",x"00",x"24",x"49",x"6d",x"92",x"b6",x"db",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"db",x"b6",x"6d",x"00",x"b6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"ed",x"c0",x"c5",x"a9",x"72",x"57",x"37",x"12",x"09",x"00",x"92",x"fa",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"e8",x"a4",x"d6",x"b7",x"00",x"00",x"00",x"b6",x"f5",x"ec",x"f0",x"f0",x"ec",x"ec",x"e8",x"c8",x"89",x"ff",x"45",x"00",x"6e",x"ff",x"ff",x"ff",x"fb",x"ff",x"ff",x"db",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"32",x"33",x"12",x"2d",x"40",x"25",x"29",x"20",x"40",x"20",x"00",x"00",x"00",x"00",x"00",x"6e",x"fa",x"ec",x"f0",x"f0",x"f0",x"ec",x"e8",x"e8",x"88",x"ff",x"6e",x"00",x"00",x"24",x"49",x"6d",x"6d",x"49",x"00",x"00",x"20",x"40",x"40",x"49",x"52",x"81",x"c0",x"c0",x"8e",x"5b",x"5b",x"5b",x"3b",x"5b",x"5b",x"7b",x"56",x"04",x"00",x"00",x"00",x"00",x"00",x"6e",x"fa",x"f0",x"f0",x"f0",x"ec",x"ec",x"e8",x"e4",x"84",x"db",x"fb",x"e8",x"e4",x"e4",x"c4",x"8d",x"ff",x"f0",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"a4",x"d6",x"ff",x"ed",x"e4",x"e8",x"e4",x"88",x"df",x"6d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"2d",x"57",x"5f",x"5f",x"3b",x"3b",x"7b",x"df",x"ff",x"49",x"00",x"00",x"00",x"24",x"92",x"b6",x"db",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"db",x"b6",x"6d",x"24",x"24",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"f2",x"c4",x"e0",x"e0",x"c4",x"89",x"6e",x"52",x"0e",x"05",x"01",x"d6",x"f5",x"ec",x"f0",x"f0",x"ec",x"ec",x"e8",x"e8",x"84",x"fb",x"6e",x"00",x"00",x"24",x"db",x"f1",x"f0",x"f0",x"f0",x"ec",x"ec",x"e8",x"a4",x"b2",x"db",x"00",x"00",x"00",x"92",x"db",x"ff",x"ff",x"df",x"b7",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"29",x"52",x"12",x"0d",x"40",x"20",x"09",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"b6",x"f5",x"ec",x"f0",x"ec",x"ec",x"ec",x"e8",x"c8",x"8d",x"ff",x"25",x"00",x"00",x"24",x"49",x"6d",x"6d",x"49",x"24",x"00",x"00",x"20",x"20",x"29",x"49",x"80",x"a0",x"84",x"72",x"3b",x"5b",x"5b",x"5b",x"5b",x"5b",x"7b",x"29",x"00",x"00",x"00",x"00",x"00",x"00",x"b6",x"fa",x"f0",x"f0",x"ec",x"ec",x"e8",x"e8",x"c4",x"a9",x"ff",x"f6",x"e4",x"e4",x"e8",x"a4",x"b6",x"fa",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e4",x"84",x"db",x"fb",x"e8",x"e4",x"e8",x"c4",x"89",x"df",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"09",x"32",x"7b",x"7b",x"7b",x"7b",x"7f",x"7f",x"9f",x"df",x"ff",x"b6",x"6d",x"49",x"49",x"24",x"6d",x"b6",x"db",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"49",x"00",x"6d",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"f6",x"c4",x"e0",x"e4",x"e0",x"e0",x"a0",x"80",x"45",x"25",x"05",x"25",x"fb",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"e8",x"c8",x"a9",x"ff",x"25",x"00",x"00",x"49",x"fb",x"f0",x"f0",x"f0",x"f0",x"ec",x"e8",x"e8",x"84",x"d6",x"b7",x"25",x"00",x"00",x"00",x"49",x"72",x"92",x"6e",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"29",x"0a",x"05",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"db",x"f1",x"f0",x"f0",x"ec",x"ec",x"ec",x"e8",x"a4",x"b2",x"db",x"00",x"00",x"00",x"24",x"49",x"49",x"6d",x"49",x"24",x"00",x"00",x"00",x"00",x"09",x"20",x"80",x"80",x"69",x"57",x"5b",x"3b",x"5b",x"5b",x"5b",x"5b",x"52",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"db",x"f5",x"f0",x"f0",x"ec",x"ec",x"e8",x"e8",x"a4",x"ad",x"ff",x"f1",x"e4",x"e4",x"e4",x"84",x"db",x"fa",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e4",x"88",x"ff",x"f6",x"e8",x"e4",x"e8",x"a4",x"b2",x"db",x"00",x"00",x"00",x"00",x"00",x"04",x"2e",x"5b",x"7f",x"7b",x"97",x"92",x"b7",x"df",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"24",x"6d",x"92",x"db",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"49",x"00",x"24",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"c9",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"60",x"20",x"00",x"4e",x"fb",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"e8",x"c4",x"ad",x"db",x"00",x"00",x"00",x"6e",x"fa",x"ec",x"f0",x"f0",x"ec",x"ec",x"e8",x"e4",x"84",x"ff",x"92",x"92",x"29",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"b6",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"05",x"05",x"25",x"25",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"fb",x"f0",x"f0",x"ec",x"ec",x"ec",x"e8",x"e8",x"a4",x"d6",x"b7",x"00",x"00",x"00",x"04",x"24",x"49",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"05",x"20",x"60",x"60",x"4e",x"37",x"57",x"3b",x"3b",x"3b",x"5b",x"57",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"ff",x"f0",x"ec",x"f0",x"ec",x"ec",x"e8",x"e8",x"a0",x"d6",x"ff",x"ed",x"e4",x"e4",x"c4",x"89",x"fb",x"f5",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"c4",x"ad",x"ff",x"f2",x"e4",x"e8",x"e8",x"84",x"db",x"92",x"00",x"00",x"00",x"00",x"05",x"52",x"7b",x"7b",x"7b",x"77",x"ae",x"a5",x"c5",x"f6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"6d",x"00",x"6d",x"92",x"db",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"49",x"24",x"00",x"49",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"c9",x"e0",x"e4",x"e0",x"e4",x"e0",x"c0",x"a0",x"a0",x"60",x"40",x"00",x"96",x"f6",x"ec",x"ec",x"f0",x"f0",x"ec",x"ec",x"e8",x"a4",x"d6",x"96",x"00",x"00",x"00",x"b6",x"f6",x"ec",x"f0",x"ec",x"ec",x"ec",x"e8",x"c4",x"89",x"ff",x"72",x"ff",x"db",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6e",x"ff",x"db",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"92",x"b6",x"b7",x"b2",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6e",x"fa",x"ec",x"f0",x"ec",x"ec",x"e8",x"e8",x"e4",x"84",x"ff",x"6e",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"49",x"24",x"20",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"05",x"0a",x"2a",x"2e",x"57",x"3b",x"5b",x"29",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6e",x"fe",x"ec",x"ec",x"f0",x"ec",x"e8",x"e8",x"e8",x"84",x"db",x"fa",x"e8",x"e4",x"e4",x"a4",x"8e",x"ff",x"f0",x"ec",x"ec",x"ec",x"e8",x"e8",x"e4",x"a0",x"b6",x"ff",x"ed",x"e4",x"e8",x"c4",x"8d",x"df",x"69",x"00",x"00",x"00",x"2e",x"5b",x"7f",x"7b",x"97",x"b2",x"a9",x"c0",x"e0",x"c0",x"c9",x"f6",x"ff",x"ff",x"ff",x"ff",x"ff",x"b6",x"00",x"24",x"6d",x"92",x"db",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"db",x"db",x"92",x"6d",x"24",x"00",x"00",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"b2",x"a5",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"80",x"60",x"20",x"00",x"d7",x"f5",x"ec",x"ec",x"f0",x"ec",x"ec",x"e8",x"e8",x"84",x"fb",x"6e",x"00",x"00",x"04",x"db",x"f1",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"a4",x"b2",x"db",x"96",x"f6",x"f6",x"db",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"b2",x"f6",x"f6",x"d7",x"45",x"00",x"00",x"00",x"25",x"b6",x"fb",x"ff",x"fa",x"fe",x"fb",x"fb",x"6e",x"00",x"00",x"00",x"00",x"00",x"00",x"b6",x"f5",x"ec",x"f0",x"ec",x"ec",x"e8",x"e8",x"c4",x"a9",x"df",x"6e",x"45",x"24",x"00",x"00",x"00",x"24",x"25",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"45",x"4d",x"4e",x"25",x"05",x"0a",x"77",x"52",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"b6",x"fa",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"c4",x"89",x"ff",x"f2",x"e4",x"e4",x"e4",x"84",x"d6",x"fa",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e4",x"84",x"db",x"fa",x"e8",x"e4",x"e8",x"a0",x"b2",x"df",x"25",x"00",x"05",x"56",x"7f",x"5b",x"7b",x"96",x"a9",x"c5",x"c4",x"e4",x"e0",x"e0",x"c0",x"c9",x"ff",x"ff",x"ff",x"ff",x"ff",x"6d",x"00",x"24",x"49",x"92",x"db",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"24",x"00",x"00",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"96",x"8d",x"c9",x"c4",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"40",x"20",x"44",x"fb",x"f1",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"c4",x"88",x"ff",x"25",x"00",x"00",x"49",x"fb",x"f0",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"a4",x"db",x"b7",x"db",x"f1",x"ec",x"fa",x"db",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"db",x"ed",x"cc",x"fa",x"fb",x"49",x"00",x"29",x"fb",x"ff",x"f5",x"d0",x"f0",x"d4",x"d0",x"f5",x"fb",x"45",x"00",x"00",x"00",x"00",x"24",x"db",x"f1",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"a4",x"d1",x"ff",x"ff",x"ff",x"fb",x"b2",x"20",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"6d",x"db",x"ff",x"ff",x"ff",x"ff",x"d7",x"29",x"25",x"00",x"00",x"00",x"00",x"24",x"6d",x"6e",x"00",x"05",x"db",x"f5",x"ec",x"f0",x"ec",x"ec",x"e8",x"e8",x"a0",x"ad",x"ff",x"ed",x"e4",x"e4",x"c4",x"64",x"ff",x"f6",x"ec",x"ec",x"ec",x"e8",x"e8",x"e4",x"e4",x"88",x"ff",x"f1",x"e4",x"e4",x"e8",x"84",x"fb",x"b7",x"00",x"2e",x"7b",x"7f",x"5b",x"76",x"8d",x"a5",x"c0",x"e0",x"e4",x"e0",x"e0",x"e0",x"c4",x"89",x"96",x"ff",x"ff",x"ff",x"ff",x"4d",x"00",x"24",x"6d",x"92",x"db",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"24",x"00",x"24",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"9f",x"7b",x"92",x"ae",x"a5",x"a4",x"c0",x"c0",x"a0",x"80",x"40",x"00",x"6d",x"fa",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"c4",x"b1",x"db",x"00",x"00",x"00",x"72",x"fa",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e4",x"84",x"db",x"92",x"fb",x"ec",x"e8",x"ec",x"fa",x"db",x"49",x"00",x"00",x"00",x"00",x"49",x"fb",x"ec",x"e8",x"f0",x"f6",x"fb",x"6e",x"d7",x"f6",x"cc",x"ec",x"ec",x"f0",x"f0",x"f0",x"cc",x"f6",x"92",x"00",x"00",x"00",x"00",x"49",x"fa",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"c4",x"d1",x"f6",x"f1",x"f1",x"f6",x"fb",x"8e",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"b2",x"fb",x"fa",x"f1",x"ed",x"ed",x"f1",x"fa",x"db",x"45",x"00",x"25",x"49",x"92",x"d6",x"ff",x"db",x"00",x"29",x"fb",x"f0",x"ec",x"ec",x"ec",x"ec",x"e8",x"e4",x"a4",x"d6",x"f6",x"e4",x"e4",x"e4",x"a0",x"92",x"ff",x"f1",x"ec",x"ec",x"ec",x"e8",x"e8",x"e4",x"c4",x"ad",x"fb",x"e8",x"e4",x"e4",x"a4",x"69",x"ff",x"6a",x"05",x"57",x"5b",x"9b",x"b2",x"a9",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c4",x"a9",x"8e",x"76",x"bb",x"ff",x"ff",x"ff",x"ff",x"92",x"00",x"24",x"6d",x"92",x"db",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"24",x"00",x"49",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"9b",x"5b",x"5b",x"7b",x"76",x"8d",x"84",x"80",x"80",x"60",x"40",x"00",x"92",x"f6",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"a4",x"d6",x"b6",x"00",x"00",x"00",x"b6",x"f5",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"c4",x"89",x"df",x"92",x"fa",x"ec",x"ec",x"e8",x"ec",x"f6",x"fb",x"69",x"00",x"00",x"00",x"6e",x"fa",x"ec",x"ec",x"ec",x"cc",x"f6",x"ff",x"f6",x"e8",x"c8",x"ec",x"ec",x"f0",x"f0",x"ec",x"ec",x"f1",x"db",x"25",x"00",x"00",x"00",x"6e",x"fa",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e4",x"e8",x"f1",x"c8",x"c8",x"c8",x"c8",x"f1",x"fb",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"92",x"ff",x"f5",x"ec",x"e8",x"e8",x"e8",x"ec",x"cc",x"f6",x"db",x"96",x"db",x"fb",x"f7",x"d2",x"fb",x"92",x"00",x"6e",x"fa",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e4",x"a4",x"f6",x"ed",x"e4",x"e4",x"e4",x"64",x"db",x"fb",x"cc",x"ec",x"ec",x"ec",x"e8",x"e8",x"e4",x"a4",x"d1",x"f2",x"e4",x"e4",x"e4",x"80",x"b2",x"db",x"25",x"2a",x"7b",x"96",x"a9",x"c4",x"e0",x"e0",x"e4",x"e4",x"e4",x"c4",x"a5",x"92",x"76",x"7b",x"5b",x"9b",x"ff",x"ff",x"ff",x"ff",x"db",x"00",x"24",x"49",x"b6",x"db",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"6d",x"24",x"00",x"92",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"9b",x"5b",x"5b",x"5b",x"7b",x"7b",x"72",x"69",x"60",x"40",x"20",x"00",x"db",x"f1",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e4",x"84",x"ff",x"6e",x"00",x"00",x"00",x"db",x"f1",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"c4",x"b2",x"db",x"b7",x"f6",x"ec",x"ec",x"ec",x"e8",x"cc",x"f6",x"fb",x"69",x"00",x"00",x"b7",x"f6",x"ec",x"ec",x"ec",x"e8",x"cc",x"f1",x"cc",x"e4",x"e8",x"e8",x"ec",x"ec",x"f0",x"ec",x"ec",x"cc",x"fb",x"49",x"00",x"00",x"00",x"b6",x"f5",x"ec",x"ec",x"ec",x"e8",x"e8",x"e4",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"ec",x"c8",x"f6",x"92",x"00",x"00",x"00",x"00",x"00",x"00",x"6e",x"ff",x"f1",x"e8",x"e8",x"e8",x"e4",x"e8",x"e8",x"ec",x"f1",x"fa",x"fa",x"f6",x"ed",x"c8",x"88",x"ff",x"6d",x"00",x"b6",x"f5",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e4",x"c8",x"ed",x"e4",x"e4",x"e4",x"a0",x"8d",x"ff",x"f6",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e4",x"c8",x"f1",x"e8",x"e4",x"e4",x"c4",x"84",x"ff",x"92",x"00",x"4e",x"ae",x"c9",x"c4",x"e0",x"e0",x"e0",x"e0",x"c0",x"a5",x"8e",x"97",x"7b",x"5b",x"3b",x"3b",x"9f",x"ff",x"fb",x"ed",x"f6",x"ff",x"48",x"04",x"6d",x"b6",x"db",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"24",x"00",x"db",x"ff",x"ff",x"ff",x"fb",x"fb",x"ff",x"ff",x"ff",x"9f",x"3b",x"5b",x"5b",x"5b",x"5b",x"57",x"52",x"49",x"20",x"00",x"49",x"fb",x"f0",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"c4",x"8d",x"ff",x"25",x"00",x"00",x"49",x"fb",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e4",x"a4",x"db",x"b7",x"d7",x"f1",x"e8",x"ec",x"ec",x"ec",x"e8",x"c8",x"d2",x"ff",x"25",x"00",x"d6",x"f1",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"c8",x"e8",x"e8",x"e8",x"ec",x"ec",x"ec",x"ec",x"ec",x"c8",x"da",x"4a",x"00",x"00",x"24",x"fb",x"f1",x"ec",x"ec",x"ec",x"e8",x"e8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"ec",x"e8",x"e8",x"d1",x"b7",x"00",x"00",x"00",x"00",x"00",x"24",x"fb",x"f5",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"ec",x"ec",x"f0",x"f0",x"e8",x"e4",x"c4",x"89",x"ff",x"25",x"20",x"fb",x"f1",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e4",x"e8",x"e8",x"e4",x"e4",x"c4",x"64",x"db",x"ff",x"f6",x"e8",x"ec",x"ec",x"e8",x"e8",x"e8",x"e4",x"e8",x"e8",x"e4",x"e4",x"e4",x"84",x"b2",x"ff",x"25",x"00",x"85",x"c5",x"e0",x"e0",x"e4",x"c0",x"a0",x"a5",x"ad",x"96",x"7b",x"5b",x"5b",x"5b",x"3b",x"3b",x"9f",x"ff",x"e9",x"e0",x"c9",x"fb",x"8d",x"00",x"6d",x"b6",x"db",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"db",x"db",x"92",x"49",x"00",x"24",x"fb",x"ff",x"ff",x"f6",x"c9",x"f2",x"ff",x"ff",x"ff",x"bf",x"5f",x"5b",x"3b",x"5b",x"3b",x"37",x"12",x"2e",x"09",x"00",x"6e",x"f6",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"c4",x"b1",x"fb",x"20",x"00",x"00",x"92",x"fa",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e4",x"84",x"fb",x"92",x"fb",x"cd",x"e8",x"ec",x"ec",x"ec",x"e8",x"c8",x"88",x"ff",x"49",x"25",x"fb",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e4",x"e4",x"a4",x"c4",x"e8",x"ec",x"ec",x"ec",x"ec",x"e8",x"c8",x"d6",x"6e",x"00",x"00",x"49",x"fb",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e4",x"e4",x"c4",x"c4",x"e8",x"e8",x"ec",x"ec",x"e8",x"c8",x"fb",x"24",x"00",x"00",x"00",x"00",x"b7",x"fa",x"ec",x"e8",x"e8",x"e4",x"c4",x"a4",x"c4",x"e8",x"e8",x"e8",x"ec",x"e8",x"e8",x"e8",x"a4",x"b2",x"db",x"00",x"49",x"fb",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e4",x"e8",x"e4",x"e4",x"e4",x"e4",x"80",x"8d",x"ff",x"ff",x"f1",x"e8",x"e8",x"ec",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"64",x"fb",x"bb",x"20",x"60",x"c0",x"e0",x"e0",x"e0",x"e0",x"a5",x"ad",x"b6",x"9b",x"5b",x"5b",x"5b",x"5b",x"5b",x"5f",x"7b",x"bb",x"cd",x"c4",x"e4",x"c4",x"a9",x"8d",x"24",x"6d",x"b6",x"db",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"db",x"ba",x"92",x"49",x"00",x"49",x"ff",x"ff",x"f2",x"e5",x"e0",x"c4",x"f2",x"ff",x"ff",x"9f",x"5b",x"5b",x"5b",x"5b",x"37",x"37",x"33",x"0e",x"09",x"00",x"b2",x"f5",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e4",x"a4",x"d6",x"b6",x"00",x"00",x"00",x"b6",x"f1",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e4",x"89",x"ff",x"92",x"fa",x"ec",x"ec",x"e8",x"ec",x"ec",x"e8",x"c4",x"8d",x"ff",x"25",x"6e",x"f6",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"80",x"64",x"ad",x"e8",x"e8",x"ec",x"ec",x"ec",x"e8",x"c4",x"d6",x"72",x"00",x"00",x"92",x"f6",x"ec",x"ec",x"ec",x"e8",x"e8",x"e4",x"e4",x"80",x"60",x"a4",x"e8",x"e8",x"e8",x"e8",x"e8",x"c8",x"db",x"49",x"00",x"00",x"00",x"6e",x"fa",x"f0",x"ec",x"e8",x"e8",x"e4",x"60",x"64",x"a8",x"e8",x"e8",x"ec",x"e8",x"e8",x"e8",x"e8",x"84",x"db",x"b6",x"00",x"6e",x"f6",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"a4",x"64",x"da",x"ff",x"fb",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"c4",x"60",x"b2",x"ff",x"4d",x"20",x"a0",x"e0",x"e0",x"c0",x"c5",x"ad",x"92",x"7b",x"7b",x"5b",x"5b",x"5b",x"5b",x"7b",x"7b",x"7b",x"96",x"ad",x"c4",x"e0",x"c4",x"a4",x"60",x"20",x"24",x"6d",x"b6",x"db",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"49",x"00",x"92",x"ff",x"d2",x"c5",x"e0",x"e0",x"e4",x"c9",x"f6",x"ff",x"9f",x"5b",x"5b",x"5b",x"5b",x"3b",x"37",x"32",x"0e",x"05",x"01",x"db",x"f1",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"e4",x"84",x"fb",x"6d",x"00",x"00",x"24",x"fb",x"f1",x"e8",x"ec",x"ec",x"e8",x"e8",x"e8",x"a4",x"b1",x"db",x"b6",x"f6",x"e8",x"ec",x"ec",x"ec",x"e8",x"e8",x"a4",x"b1",x"db",x"01",x"b3",x"f6",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e4",x"84",x"d6",x"fa",x"ec",x"e8",x"ec",x"ec",x"ec",x"e8",x"c4",x"d6",x"72",x"00",x"00",x"b7",x"f5",x"ec",x"ec",x"ec",x"e8",x"e8",x"e4",x"e4",x"84",x"d6",x"f6",x"e8",x"e8",x"e8",x"e8",x"e8",x"c8",x"fb",x"49",x"00",x"00",x"24",x"db",x"f5",x"ec",x"ec",x"e8",x"e8",x"c4",x"89",x"d6",x"f1",x"e8",x"e8",x"e8",x"ec",x"e8",x"e8",x"e4",x"84",x"ff",x"6d",x"00",x"b7",x"f5",x"e8",x"ec",x"ec",x"ec",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"c4",x"60",x"b2",x"ff",x"ff",x"f6",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e8",x"80",x"89",x"ff",x"b6",x"00",x"60",x"e0",x"e0",x"c5",x"89",x"b2",x"97",x"7b",x"5b",x"5b",x"3b",x"5b",x"5b",x"5b",x"7b",x"97",x"ae",x"a9",x"c5",x"c4",x"80",x"40",x"40",x"20",x"00",x"29",x"92",x"b6",x"db",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"db",x"db",x"92",x"49",x"20",x"d6",x"f2",x"c4",x"e0",x"e4",x"e0",x"e0",x"e0",x"c9",x"fb",x"bf",x"5b",x"5f",x"3b",x"3b",x"3b",x"37",x"12",x"09",x"00",x"25",x"fb",x"ec",x"e8",x"ec",x"ec",x"e8",x"e8",x"e8",x"c4",x"a9",x"ff",x"49",x"00",x"00",x"49",x"fb",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"84",x"da",x"b7",x"db",x"f1",x"e8",x"ec",x"ec",x"ec",x"e8",x"e4",x"a4",x"da",x"92",x"01",x"db",x"f1",x"e8",x"ec",x"ec",x"e8",x"e8",x"e4",x"c4",x"ad",x"ff",x"ff",x"ec",x"e8",x"ec",x"e8",x"e8",x"e8",x"c4",x"d6",x"92",x"00",x"04",x"fb",x"f1",x"e8",x"ec",x"e8",x"e8",x"e8",x"e4",x"c0",x"ad",x"ff",x"fb",x"ec",x"e8",x"e8",x"e8",x"e8",x"a4",x"fb",x"6d",x"00",x"00",x"6e",x"fb",x"ec",x"ec",x"e8",x"e8",x"e4",x"a4",x"d6",x"ff",x"f6",x"e8",x"e8",x"ec",x"ec",x"e8",x"e8",x"c4",x"89",x"ff",x"24",x"00",x"fb",x"f1",x"e8",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"60",x"89",x"ff",x"db",x"db",x"f6",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"c4",x"64",x"db",x"ff",x"49",x"20",x"80",x"c0",x"a9",x"92",x"97",x"7b",x"5b",x"5b",x"5f",x"3f",x"5b",x"9b",x"9b",x"76",x"8e",x"a9",x"c5",x"a4",x"80",x"60",x"20",x"00",x"00",x"00",x"24",x"69",x"92",x"b6",x"db",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"49",x"24",x"ae",x"a4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c4",x"c9",x"b7",x"7b",x"5b",x"5b",x"3b",x"37",x"13",x"0e",x"09",x"00",x"6e",x"fa",x"e8",x"e8",x"ec",x"ec",x"e8",x"e8",x"e4",x"a4",x"d2",x"db",x"00",x"00",x"00",x"72",x"f6",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"88",x"ff",x"92",x"fb",x"ec",x"e8",x"ec",x"ec",x"e8",x"e8",x"e4",x"a8",x"fb",x"4a",x"25",x"fb",x"ec",x"e8",x"ec",x"ec",x"e8",x"e8",x"e4",x"a4",x"d2",x"ff",x"fa",x"e8",x"e8",x"ec",x"e8",x"e8",x"e4",x"a4",x"d6",x"6e",x"00",x"49",x"fb",x"ec",x"e8",x"ec",x"e8",x"e8",x"e4",x"e4",x"a0",x"d6",x"ff",x"fa",x"e8",x"e8",x"e8",x"e8",x"e8",x"a4",x"fb",x"49",x"00",x"04",x"db",x"f5",x"ec",x"ec",x"e8",x"e8",x"e4",x"84",x"db",x"ff",x"f6",x"e8",x"e8",x"ec",x"ec",x"e8",x"e4",x"a4",x"b2",x"db",x"00",x"49",x"fb",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"80",x"64",x"db",x"df",x"4e",x"db",x"f1",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"a4",x"60",x"b6",x"ff",x"72",x"00",x"20",x"89",x"92",x"76",x"7b",x"7b",x"5b",x"3b",x"5b",x"5b",x"5b",x"97",x"92",x"8d",x"a9",x"a4",x"a4",x"60",x"40",x"20",x"00",x"00",x"00",x"04",x"24",x"49",x"6d",x"b2",x"db",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"49",x"20",x"44",x"80",x"c4",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c9",x"92",x"76",x"77",x"57",x"37",x"33",x"0e",x"05",x"00",x"96",x"f6",x"e8",x"ec",x"e8",x"e8",x"e8",x"e8",x"e4",x"a4",x"db",x"b7",x"00",x"00",x"00",x"b7",x"f1",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"a0",x"8d",x"df",x"72",x"fa",x"e8",x"e8",x"ec",x"e8",x"e8",x"e8",x"c4",x"ad",x"ff",x"25",x"6e",x"fa",x"e8",x"ec",x"ec",x"e8",x"e8",x"e4",x"e4",x"84",x"db",x"ff",x"f6",x"e8",x"e8",x"ec",x"e8",x"e8",x"e4",x"a4",x"db",x"6d",x"00",x"92",x"fa",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"84",x"fb",x"ff",x"f6",x"c8",x"e8",x"e8",x"e8",x"e8",x"a4",x"fb",x"49",x"00",x"4d",x"fb",x"ec",x"e8",x"e8",x"e8",x"e4",x"e4",x"89",x"ff",x"ff",x"d1",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"a4",x"db",x"92",x"00",x"72",x"f6",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"a0",x"60",x"d6",x"ff",x"72",x"29",x"fb",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"c0",x"60",x"91",x"ff",x"db",x"00",x"00",x"6d",x"97",x"7b",x"5b",x"5b",x"5f",x"3f",x"5b",x"7b",x"97",x"92",x"ae",x"a5",x"a4",x"80",x"60",x"20",x"00",x"00",x"00",x"00",x"04",x"24",x"29",x"49",x"6d",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"20",x"20",x"20",x"40",x"40",x"80",x"c0",x"c4",x"e4",x"e0",x"e0",x"e0",x"c5",x"a9",x"8d",x"72",x"52",x"32",x"09",x"05",x"00",x"db",x"f1",x"e8",x"ec",x"e8",x"e8",x"e8",x"e4",x"e4",x"84",x"fb",x"6e",x"00",x"00",x"24",x"fb",x"ed",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"80",x"d7",x"b7",x"96",x"f6",x"e8",x"e8",x"ec",x"e8",x"e8",x"e8",x"a4",x"b2",x"db",x"01",x"b2",x"f5",x"e8",x"ec",x"ec",x"e8",x"e8",x"e4",x"c4",x"84",x"ff",x"ff",x"f1",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"84",x"db",x"69",x"00",x"b7",x"f1",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"c4",x"89",x"ff",x"fb",x"f1",x"e8",x"e8",x"e8",x"e8",x"e4",x"a8",x"fb",x"45",x"00",x"b6",x"f6",x"e8",x"e8",x"e8",x"e8",x"e4",x"c4",x"b2",x"ff",x"fb",x"cc",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"88",x"ff",x"4d",x"00",x"b6",x"f1",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"80",x"64",x"b2",x"ff",x"b7",x"21",x"6e",x"fa",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"a0",x"60",x"8d",x"ff",x"ff",x"49",x"00",x"2d",x"77",x"5b",x"3f",x"5f",x"5b",x"5b",x"7b",x"97",x"b2",x"a9",x"a5",x"c4",x"e9",x"cd",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"48",x"49",x"49",x"6d",x"92",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"24",x"00",x"00",x"00",x"00",x"20",x"40",x"60",x"a0",x"c4",x"c4",x"e0",x"c0",x"c0",x"a0",x"85",x"65",x"29",x"05",x"00",x"29",x"fb",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"c4",x"89",x"ff",x"25",x"00",x"00",x"b2",x"f6",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"c4",x"89",x"ff",x"6e",x"b7",x"f1",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"84",x"db",x"92",x"01",x"db",x"ed",x"e8",x"ec",x"e8",x"e8",x"e8",x"e4",x"c0",x"8d",x"ff",x"fb",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"89",x"fb",x"49",x"01",x"fb",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"a4",x"b2",x"ff",x"fb",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"ad",x"db",x"25",x"25",x"fb",x"ed",x"e8",x"e8",x"e8",x"e4",x"e4",x"a0",x"d6",x"ff",x"f6",x"c8",x"e8",x"e8",x"e8",x"e8",x"e4",x"c4",x"89",x"ff",x"25",x"20",x"fb",x"ed",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"80",x"68",x"b6",x"ff",x"db",x"25",x"00",x"b6",x"f6",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"a0",x"84",x"91",x"ff",x"ff",x"6e",x"00",x"05",x"57",x"5b",x"3f",x"5b",x"7b",x"7b",x"97",x"92",x"a9",x"a5",x"a0",x"c0",x"e0",x"e9",x"d6",x"00",x"00",x"00",x"00",x"24",x"45",x"69",x"69",x"6d",x"8e",x"92",x"92",x"ba",x"db",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"49",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"20",x"40",x"60",x"a0",x"c0",x"e0",x"c0",x"a0",x"80",x"40",x"00",x"00",x"6e",x"fa",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"a0",x"d2",x"db",x"00",x"00",x"49",x"fb",x"f1",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"80",x"b6",x"ff",x"4a",x"db",x"ec",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"84",x"ff",x"49",x"25",x"fb",x"cc",x"e8",x"ec",x"e8",x"e8",x"e8",x"e4",x"a0",x"d2",x"ff",x"fa",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"c0",x"ad",x"db",x"04",x"49",x"fb",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"80",x"d6",x"ff",x"fa",x"e8",x"e8",x"e8",x"e8",x"e8",x"c0",x"b1",x"db",x"00",x"6e",x"fa",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"84",x"db",x"ff",x"f2",x"e4",x"e8",x"e8",x"e8",x"e4",x"e4",x"a0",x"d2",x"db",x"00",x"49",x"fb",x"ec",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"a4",x"89",x"db",x"ff",x"db",x"49",x"00",x"00",x"db",x"f1",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"c4",x"64",x"b2",x"ff",x"ff",x"8e",x"00",x"05",x"33",x"5b",x"5f",x"7f",x"7b",x"92",x"b2",x"a9",x"a4",x"a4",x"a5",x"84",x"c4",x"e4",x"c4",x"fb",x"49",x"00",x"00",x"04",x"24",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b2",x"71",x"4d",x"49",x"45",x"24",x"24",x"00",x"00",x"00",x"00",x"20",x"40",x"60",x"a0",x"a0",x"a0",x"80",x"40",x"20",x"00",x"b6",x"f2",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"a4",x"fb",x"b2",x"00",x"24",x"b7",x"f6",x"e8",x"e4",x"e8",x"e4",x"e4",x"e4",x"c0",x"68",x"ff",x"97",x"49",x"fa",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"c0",x"a9",x"df",x"25",x"6e",x"fa",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"a4",x"db",x"ff",x"f2",x"e4",x"e4",x"e8",x"e8",x"e4",x"e8",x"a0",x"b2",x"db",x"00",x"92",x"f6",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"84",x"fb",x"ff",x"f1",x"e4",x"e8",x"e8",x"e8",x"e4",x"a0",x"d6",x"b7",x"01",x"b7",x"f1",x"e8",x"e8",x"e8",x"e8",x"e4",x"c4",x"89",x"ff",x"ff",x"ed",x"e4",x"e8",x"e8",x"e8",x"e4",x"e4",x"80",x"fb",x"92",x"00",x"92",x"f6",x"c8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"84",x"db",x"ff",x"db",x"49",x"00",x"00",x"49",x"fb",x"ec",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"a0",x"b2",x"ff",x"ff",x"92",x"00",x"00",x"2e",x"7b",x"5b",x"7b",x"96",x"b2",x"a9",x"a4",x"80",x"84",x"ad",x"b2",x"d6",x"cd",x"e4",x"c4",x"f6",x"6e",x"00",x"00",x"24",x"49",x"6d",x"72",x"96",x"b6",x"b6",x"ba",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"6d",x"6d",x"49",x"49",x"44",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"20",x"40",x"40",x"40",x"40",x"20",x"00",x"db",x"ed",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"84",x"fb",x"6e",x"05",x"b2",x"fa",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"84",x"b6",x"ff",x"25",x"92",x"f6",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"a0",x"d2",x"bb",x"01",x"96",x"f1",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"84",x"ff",x"ff",x"ed",x"e4",x"e8",x"e8",x"e4",x"e4",x"e4",x"80",x"da",x"92",x"00",x"b6",x"f1",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"c4",x"8d",x"ff",x"fb",x"ed",x"e4",x"e8",x"e8",x"e4",x"e4",x"a4",x"fb",x"6e",x"25",x"fb",x"ec",x"e8",x"e8",x"e8",x"e4",x"e4",x"a0",x"b1",x"ff",x"fb",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"c4",x"84",x"ff",x"49",x"00",x"b7",x"f1",x"e4",x"e8",x"e8",x"e8",x"e8",x"e4",x"c4",x"89",x"ff",x"bb",x"49",x"00",x"00",x"00",x"6e",x"f6",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"84",x"fb",x"db",x"6e",x"00",x"00",x"09",x"57",x"97",x"96",x"8e",x"a5",x"c5",x"c0",x"80",x"64",x"b2",x"ff",x"ff",x"ff",x"fb",x"e4",x"c4",x"d2",x"92",x"00",x"24",x"49",x"6d",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"b6",x"92",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"25",x"fb",x"cc",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"c4",x"89",x"ff",x"49",x"92",x"fb",x"ed",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"80",x"69",x"ff",x"96",x"01",x"db",x"f1",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"80",x"fa",x"92",x"01",x"db",x"ed",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"c0",x"a9",x"ff",x"fb",x"ec",x"e4",x"e8",x"e8",x"e4",x"e4",x"c4",x"84",x"ff",x"4d",x"05",x"fb",x"ed",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"a0",x"b2",x"ff",x"fb",x"e8",x"e4",x"e8",x"e4",x"e4",x"e4",x"a4",x"fb",x"49",x"4a",x"fa",x"c8",x"e8",x"e8",x"e8",x"e4",x"e4",x"a0",x"d6",x"df",x"f6",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"c4",x"ad",x"db",x"25",x"00",x"db",x"ed",x"e4",x"e8",x"e8",x"e8",x"e4",x"e4",x"a0",x"d2",x"df",x"25",x"00",x"00",x"00",x"00",x"b6",x"f6",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"c4",x"a8",x"ff",x"6d",x"00",x"00",x"24",x"72",x"92",x"ad",x"a9",x"c4",x"e4",x"e4",x"c4",x"64",x"d6",x"ff",x"ff",x"db",x"bb",x"fb",x"e8",x"c0",x"d2",x"96",x"00",x"24",x"49",x"6e",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"49",x"45",x"24",x"04",x"00",x"00",x"00",x"00",x"00",x"6d",x"f6",x"c8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"a0",x"b2",x"ff",x"db",x"fa",x"e9",x"e4",x"e8",x"e4",x"e4",x"e4",x"e4",x"a0",x"64",x"db",x"fb",x"25",x"25",x"fb",x"ec",x"e4",x"e8",x"e4",x"e4",x"e4",x"e4",x"84",x"ff",x"4a",x"25",x"fb",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"a0",x"b2",x"ff",x"fa",x"c8",x"e4",x"e8",x"e8",x"e4",x"e4",x"c0",x"ad",x"ff",x"25",x"29",x"fb",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"a0",x"da",x"ff",x"f6",x"c8",x"e4",x"e8",x"e4",x"e4",x"c0",x"a9",x"ff",x"25",x"92",x"f6",x"c8",x"e8",x"e8",x"e8",x"e4",x"e4",x"a4",x"fb",x"df",x"f2",x"e4",x"e8",x"e8",x"e8",x"e4",x"e4",x"a0",x"d2",x"db",x"00",x"49",x"fb",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"a4",x"d6",x"96",x"00",x"00",x"00",x"00",x"00",x"db",x"ed",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"c0",x"ad",x"db",x"20",x"00",x"00",x"44",x"a9",x"85",x"64",x"a9",x"f1",x"e8",x"c4",x"64",x"b2",x"ff",x"db",x"72",x"24",x"29",x"db",x"e8",x"c0",x"b2",x"b6",x"00",x"24",x"49",x"92",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"69",x"49",x"45",x"24",x"00",x"00",x"00",x"00",x"b6",x"f6",x"c4",x"e8",x"e8",x"e8",x"e4",x"e4",x"e0",x"a0",x"d6",x"ff",x"f6",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a4",x"40",x"b2",x"ff",x"92",x"00",x"49",x"fb",x"c8",x"e4",x"e8",x"e4",x"e4",x"e4",x"c0",x"8d",x"ff",x"25",x"6e",x"f6",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"a0",x"db",x"ff",x"f2",x"c4",x"e8",x"e8",x"e4",x"e4",x"e4",x"a0",x"b2",x"db",x"00",x"72",x"f6",x"e4",x"e8",x"e8",x"e8",x"e4",x"e4",x"c0",x"a4",x"ff",x"ff",x"f2",x"e4",x"e4",x"e8",x"e4",x"e4",x"c0",x"b2",x"db",x"25",x"d7",x"ed",x"e4",x"e8",x"e8",x"e4",x"e4",x"c4",x"a9",x"ff",x"ff",x"cd",x"e4",x"e8",x"e8",x"e4",x"e4",x"e4",x"80",x"d6",x"92",x"00",x"6e",x"f6",x"e4",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"84",x"fb",x"6e",x"00",x"00",x"00",x"00",x"29",x"fb",x"c8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"a0",x"d6",x"b7",x"00",x"00",x"00",x"44",x"60",x"40",x"00",x"d2",x"f2",x"e4",x"80",x"69",x"ff",x"db",x"49",x"00",x"00",x"04",x"db",x"e8",x"c0",x"d6",x"b6",x"00",x"24",x"6d",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"49",x"44",x"20",x"00",x"00",x"00",x"fb",x"ed",x"e4",x"e8",x"e8",x"e4",x"e4",x"e4",x"e0",x"c4",x"fa",x"ed",x"e4",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"64",x"b6",x"ff",x"d7",x"00",x"00",x"92",x"f2",x"e4",x"e4",x"e8",x"e4",x"e4",x"e4",x"a0",x"d6",x"db",x"01",x"b7",x"f1",x"e4",x"e8",x"e8",x"e4",x"e4",x"e4",x"c0",x"84",x"ff",x"ff",x"ed",x"e4",x"e8",x"e4",x"e4",x"e4",x"e4",x"80",x"db",x"92",x"00",x"b7",x"f1",x"e4",x"e8",x"e8",x"e4",x"e4",x"e4",x"c0",x"a9",x"ff",x"fb",x"ed",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"d6",x"96",x"25",x"fb",x"e8",x"e4",x"e4",x"e8",x"e4",x"e4",x"a0",x"b2",x"ff",x"fb",x"c8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a4",x"ff",x"49",x"00",x"b7",x"f1",x"e4",x"e8",x"e8",x"e4",x"e4",x"e4",x"c0",x"89",x"ff",x"25",x"00",x"00",x"00",x"00",x"6e",x"fa",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"84",x"fb",x"72",x"00",x"00",x"00",x"00",x"00",x"00",x"6e",x"f6",x"e4",x"e0",x"64",x"db",x"ff",x"49",x"00",x"00",x"00",x"25",x"fb",x"e4",x"a0",x"da",x"92",x"00",x"28",x"6d",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"92",x"72",x"6d",x"49",x"24",x"00",x"00",x"29",x"fb",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"ed",x"e4",x"e0",x"e0",x"e4",x"e4",x"e0",x"c0",x"80",x"60",x"b2",x"ff",x"db",x"25",x"00",x"00",x"d7",x"f1",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"80",x"fb",x"92",x"01",x"db",x"ed",x"e4",x"e8",x"e8",x"e4",x"e4",x"e4",x"c0",x"ad",x"ff",x"fb",x"e8",x"e4",x"e8",x"e4",x"e4",x"e4",x"e4",x"84",x"df",x"49",x"25",x"fb",x"e8",x"e4",x"e8",x"e8",x"e4",x"e4",x"e4",x"a0",x"b2",x"ff",x"fa",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"84",x"ff",x"4e",x"4e",x"f6",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"80",x"d6",x"ff",x"f6",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"ad",x"ff",x"25",x"25",x"fb",x"ed",x"e4",x"e8",x"e8",x"e4",x"e4",x"e4",x"a0",x"b2",x"db",x"00",x"00",x"00",x"00",x"00",x"b6",x"f1",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"c0",x"89",x"ff",x"49",x"00",x"00",x"00",x"00",x"00",x"25",x"db",x"cd",x"e0",x"80",x"91",x"ff",x"4e",x"00",x"00",x"00",x"00",x"49",x"f6",x"e4",x"a4",x"db",x"6d",x"00",x"49",x"6d",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"96",x"92",x"6d",x"49",x"24",x"00",x"00",x"6e",x"f6",x"e8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"e0",x"e4",x"e4",x"c4",x"c0",x"a0",x"40",x"69",x"db",x"ff",x"fb",x"49",x"00",x"00",x"25",x"fa",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"84",x"ff",x"49",x"29",x"fb",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"b2",x"ff",x"f6",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"ad",x"df",x"25",x"49",x"fa",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a4",x"db",x"ff",x"f6",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"88",x"ff",x"25",x"92",x"f2",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"84",x"df",x"ff",x"f1",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"b2",x"db",x"00",x"49",x"fb",x"e8",x"e4",x"e8",x"e4",x"e4",x"e4",x"e4",x"a0",x"d7",x"96",x"00",x"00",x"00",x"00",x"24",x"db",x"ed",x"e4",x"e8",x"e4",x"e4",x"e4",x"e4",x"a0",x"ad",x"db",x"00",x"00",x"00",x"00",x"00",x"00",x"b2",x"f2",x"e4",x"c4",x"64",x"fb",x"d7",x"00",x"00",x"00",x"00",x"00",x"92",x"f2",x"c0",x"84",x"fb",x"29",x"00",x"49",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"d6",x"b6",x"92",x"49",x"24",x"00",x"00",x"b3",x"f2",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"e0",x"e0",x"e0",x"c4",x"c0",x"80",x"60",x"44",x"92",x"df",x"ff",x"ff",x"49",x"00",x"00",x"00",x"6e",x"fa",x"e8",x"e4",x"e8",x"e4",x"e4",x"e4",x"c0",x"89",x"ff",x"01",x"6e",x"f6",x"e4",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"d6",x"ff",x"f2",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"b2",x"db",x"00",x"92",x"f6",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"84",x"ff",x"df",x"f1",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"ad",x"db",x"25",x"db",x"ed",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"89",x"ff",x"ff",x"ed",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"80",x"da",x"96",x"00",x"6e",x"f6",x"e4",x"e4",x"e8",x"e4",x"e4",x"e4",x"e0",x"84",x"ff",x"72",x"00",x"00",x"00",x"00",x"49",x"fb",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"d6",x"b7",x"00",x"00",x"00",x"00",x"00",x"4d",x"fb",x"e8",x"e0",x"80",x"91",x"ff",x"6a",x"00",x"00",x"00",x"00",x"00",x"b7",x"ed",x"c0",x"89",x"ff",x"25",x"00",x"49",x"92",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"92",x"49",x"24",x"00",x"00",x"db",x"ed",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"a0",x"60",x"60",x"60",x"40",x"64",x"89",x"b6",x"ff",x"ff",x"ff",x"d7",x"25",x"00",x"00",x"00",x"00",x"b6",x"f1",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"a0",x"b6",x"db",x"01",x"b7",x"f1",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"84",x"ff",x"ff",x"ed",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"80",x"db",x"92",x"00",x"d7",x"ed",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"c0",x"8d",x"ff",x"fb",x"ed",x"e0",x"e4",x"e4",x"e4",x"e0",x"c0",x"d1",x"db",x"92",x"fb",x"e8",x"e4",x"e4",x"e4",x"e4",x"e0",x"a0",x"b2",x"ff",x"fb",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"84",x"fb",x"6a",x"00",x"b7",x"ed",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"89",x"ff",x"25",x"00",x"00",x"00",x"00",x"8e",x"f6",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"84",x"fb",x"72",x"00",x"00",x"00",x"00",x"20",x"db",x"ed",x"e4",x"e0",x"64",x"fb",x"b7",x"00",x"00",x"00",x"00",x"00",x"49",x"f6",x"e4",x"a0",x"b2",x"db",x"00",x"24",x"49",x"92",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"49",x"24",x"00",x"49",x"fb",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"c0",x"84",x"89",x"ad",x"ad",x"b2",x"da",x"fb",x"ff",x"ff",x"ff",x"92",x"24",x"00",x"00",x"00",x"00",x"00",x"d7",x"ed",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"d7",x"92",x"01",x"db",x"ed",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"89",x"ff",x"ff",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"a4",x"ff",x"69",x"25",x"fb",x"ed",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"a0",x"b2",x"ff",x"fb",x"c4",x"e0",x"e4",x"e4",x"e4",x"e4",x"c0",x"ed",x"fb",x"fb",x"f2",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"a0",x"d6",x"ff",x"f6",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"ad",x"fb",x"25",x"05",x"fb",x"ed",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"b2",x"db",x"00",x"00",x"00",x"00",x"00",x"db",x"f1",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"a9",x"ff",x"49",x"00",x"00",x"00",x"00",x"92",x"f6",x"c4",x"e0",x"a0",x"8d",x"ff",x"6d",x"00",x"00",x"00",x"00",x"00",x"92",x"f2",x"e4",x"80",x"d6",x"b6",x"00",x"24",x"6d",x"92",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"49",x"24",x"00",x"6e",x"f6",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"ad",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"b6",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"f7",x"e8",x"e0",x"e4",x"e4",x"e4",x"e4",x"e0",x"84",x"ff",x"45",x"29",x"fb",x"c8",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"a0",x"b2",x"ff",x"f6",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"ad",x"ff",x"20",x"69",x"fb",x"c8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"a4",x"db",x"ff",x"f6",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"ed",x"ed",x"c4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"a4",x"fb",x"ff",x"f2",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"d2",x"bb",x"00",x"6d",x"f7",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"db",x"b6",x"00",x"00",x"00",x"00",x"b6",x"f6",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"ad",x"db",x"00",x"00",x"00",x"00",x"6e",x"fb",x"c9",x"e0",x"c0",x"60",x"db",x"db",x"00",x"00",x"00",x"00",x"00",x"25",x"db",x"c9",x"c0",x"84",x"ff",x"6d",x"00",x"24",x"6d",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"49",x"20",x"00",x"b6",x"f1",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"a0",x"da",x"ff",x"ff",x"ff",x"db",x"96",x"6e",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6e",x"f6",x"e4",x"e0",x"e4",x"e4",x"e0",x"e0",x"c0",x"8d",x"ff",x"49",x"b6",x"f2",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"80",x"b6",x"ff",x"f1",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"b2",x"bb",x"49",x"d7",x"f2",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"88",x"ff",x"ff",x"ed",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e4",x"e4",x"e4",x"e4",x"e0",x"c0",x"a9",x"ff",x"ff",x"e9",x"e0",x"e4",x"e4",x"e4",x"e4",x"e0",x"a0",x"fb",x"96",x"49",x"fb",x"ed",x"c0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"a4",x"ff",x"6e",x"00",x"00",x"20",x"b2",x"fb",x"c9",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c0",x"d6",x"b7",x"00",x"00",x"00",x"6e",x"fb",x"ed",x"c0",x"e0",x"80",x"8d",x"ff",x"6e",x"00",x"00",x"00",x"00",x"00",x"6e",x"f6",x"c4",x"a0",x"ad",x"ff",x"24",x"00",x"49",x"91",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"6d",x"49",x"00",x"00",x"db",x"e9",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"84",x"df",x"92",x"45",x"25",x"25",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"b2",x"ed",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"d1",x"ff",x"d6",x"f6",x"e9",x"e0",x"e0",x"e4",x"e4",x"e4",x"e0",x"e0",x"84",x"df",x"ff",x"e9",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"c4",x"f6",x"df",x"d7",x"f6",x"c8",x"e0",x"e4",x"e4",x"e4",x"e4",x"e0",x"c0",x"ad",x"ff",x"fb",x"e9",x"e0",x"e4",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"a0",x"b2",x"df",x"fb",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"c4",x"fb",x"db",x"f7",x"f2",x"e4",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"c4",x"ff",x"29",x"00",x"69",x"d6",x"f6",x"c9",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"c4",x"fa",x"72",x"00",x"45",x"b2",x"f7",x"ed",x"e0",x"e0",x"c0",x"64",x"db",x"df",x"25",x"00",x"00",x"00",x"00",x"25",x"d6",x"e9",x"e0",x"80",x"d6",x"bb",x"00",x"00",x"49",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"6d",x"24",x"00",x"49",x"fb",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"c0",x"a9",x"ff",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"d7",x"e9",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e9",x"fb",x"f2",x"e9",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e0",x"c0",x"89",x"ff",x"fb",x"e4",x"e0",x"e4",x"e4",x"e4",x"e4",x"e0",x"e4",x"f1",x"fb",x"f2",x"e5",x"e0",x"e0",x"e4",x"e4",x"e4",x"e0",x"e0",x"c0",x"b2",x"ff",x"fa",x"e4",x"e0",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e0",x"e4",x"e4",x"e0",x"e0",x"a0",x"d6",x"ff",x"f6",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"c4",x"f6",x"f6",x"ed",x"c4",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"c4",x"fb",x"b6",x"b2",x"f6",x"f6",x"c9",x"c0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"c4",x"f6",x"db",x"92",x"d7",x"f6",x"ed",x"e0",x"e0",x"e4",x"80",x"8d",x"ff",x"92",x"00",x"00",x"00",x"00",x"00",x"92",x"f6",x"e0",x"c0",x"84",x"ff",x"6e",x"00",x"24",x"49",x"92",x"da",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"92",x"49",x"24",x"00",x"6e",x"f6",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"a0",x"d2",x"db",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"f7",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c8",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"b2",x"ff",x"f6",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e0",x"e0",x"e4",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"c0",x"d6",x"ff",x"f2",x"e0",x"e0",x"e0",x"e4",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e0",x"e0",x"a4",x"fb",x"ff",x"ed",x"e0",x"e0",x"e4",x"e4",x"e0",x"e4",x"e0",x"e0",x"e8",x"e9",x"c0",x"c0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e0",x"e4",x"f1",x"f6",x"f6",x"ed",x"c4",x"c0",x"e0",x"e0",x"e4",x"e0",x"e4",x"e4",x"e4",x"e0",x"e0",x"e4",x"ed",x"f6",x"f2",x"f2",x"c9",x"e0",x"e0",x"e0",x"a0",x"64",x"db",x"db",x"24",x"00",x"00",x"00",x"00",x"25",x"f7",x"e9",x"c0",x"80",x"b2",x"ff",x"25",x"00",x"24",x"6d",x"92",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"49",x"24",x"00",x"b7",x"ed",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"a0",x"db",x"96",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"f6",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"80",x"d6",x"ff",x"f2",x"e0",x"e4",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c4",x"fb",x"ff",x"c9",x"e0",x"e0",x"e0",x"e0",x"80",x"a4",x"c0",x"c0",x"c0",x"a0",x"a0",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c4",x"ff",x"fb",x"e4",x"e0",x"e0",x"e4",x"e4",x"e0",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e0",x"e0",x"e4",x"e0",x"e4",x"e4",x"e9",x"e4",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"c0",x"60",x"b6",x"ff",x"6e",x"00",x"00",x"00",x"00",x"00",x"b2",x"f2",x"e0",x"c0",x"84",x"db",x"b7",x"00",x"00",x"48",x"6d",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"6d",x"49",x"00",x"00",x"db",x"c9",x"e0",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"84",x"ff",x"6d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"69",x"f2",x"a0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"84",x"db",x"fb",x"ed",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c4",x"f6",x"f6",x"c4",x"e0",x"e0",x"e0",x"a0",x"89",x"d2",x"84",x"80",x"60",x"64",x"a9",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c4",x"fa",x"f1",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"80",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"89",x"ff",x"bb",x"00",x"00",x"00",x"00",x"00",x"4e",x"f7",x"e9",x"e0",x"80",x"8d",x"ff",x"6d",x"00",x"00",x"49",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"6d",x"24",x"00",x"49",x"f7",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"8d",x"ff",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"45",x"49",x"49",x"69",x"6e",x"6e",x"8e",x"8e",x"b6",x"d6",x"84",x"84",x"a4",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"89",x"db",x"db",x"ed",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a0",x"e0",x"e0",x"e4",x"e0",x"e0",x"e0",x"e4",x"ed",x"e9",x"e0",x"e0",x"e0",x"c0",x"60",x"b6",x"ff",x"b6",x"8d",x"8e",x"b6",x"f6",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c4",x"e9",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"a4",x"c4",x"e0",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"89",x"c9",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"80",x"69",x"db",x"ff",x"49",x"00",x"00",x"00",x"00",x"25",x"d7",x"ed",x"e0",x"c0",x"60",x"db",x"db",x"00",x"00",x"24",x"6d",x"92",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"4d",x"04",x"00",x"8e",x"f2",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"d2",x"db",x"00",x"00",x"00",x"24",x"49",x"72",x"b6",x"d7",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"d2",x"d2",x"b1",x"ad",x"ad",x"88",x"a4",x"84",x"80",x"80",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"ad",x"bb",x"bb",x"ed",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"68",x"c9",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"ad",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"60",x"89",x"d6",x"c8",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"60",x"89",x"ff",x"cd",x"c0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"80",x"65",x"db",x"ff",x"92",x"00",x"00",x"00",x"00",x"00",x"b2",x"f6",x"c0",x"e0",x"a0",x"89",x"ff",x"6e",x"00",x"00",x"49",x"6d",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"49",x"00",x"00",x"b6",x"ed",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"da",x"96",x"21",x"45",x"8e",x"b6",x"fb",x"fb",x"fb",x"f7",x"f6",x"f2",x"ed",x"ed",x"ed",x"ed",x"e9",x"e9",x"ed",x"ed",x"ed",x"f1",x"f2",x"f2",x"f2",x"f2",x"d2",x"ad",x"89",x"84",x"84",x"84",x"a0",x"a0",x"c0",x"c0",x"e0",x"a0",x"d6",x"72",x"b6",x"f1",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"68",x"da",x"f6",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"69",x"fb",x"ff",x"92",x"b7",x"db",x"db",x"bb",x"ff",x"c9",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"69",x"db",x"ff",x"d2",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"60",x"89",x"db",x"ff",x"f6",x"a4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"64",x"b6",x"ff",x"b7",x"21",x"00",x"00",x"00",x"00",x"6e",x"f6",x"e4",x"e0",x"c0",x"80",x"d7",x"db",x"24",x"00",x"24",x"49",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"6d",x"49",x"00",x"00",x"fb",x"c9",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"84",x"ff",x"b7",x"b2",x"fb",x"fb",x"f6",x"f2",x"e9",x"e5",x"e0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"e4",x"e9",x"ed",x"f2",x"f6",x"f6",x"f6",x"d6",x"b1",x"ad",x"84",x"80",x"a0",x"a0",x"84",x"fb",x"25",x"92",x"f6",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"69",x"db",x"ff",x"ff",x"a5",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"80",x"89",x"fb",x"ff",x"6e",x"00",x"00",x"49",x"49",x"24",x"db",x"f2",x"a0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"a4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"60",x"8d",x"ff",x"ff",x"ff",x"fb",x"a9",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"60",x"8d",x"ff",x"ff",x"db",x"ff",x"cd",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"60",x"69",x"da",x"ff",x"db",x"25",x"00",x"00",x"00",x"00",x"6d",x"fb",x"e9",x"e0",x"e0",x"80",x"ad",x"ff",x"6e",x"00",x"00",x"24",x"6d",x"92",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"6d",x"24",x"00",x"49",x"f6",x"a4",x"c0",x"e0",x"c0",x"e0",x"e0",x"e0",x"a0",x"a9",x"ff",x"fb",x"f6",x"f2",x"e9",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c4",x"e8",x"ed",x"f1",x"f6",x"f6",x"f6",x"d2",x"ad",x"64",x"89",x"db",x"05",x"6e",x"fb",x"a9",x"a0",x"e0",x"c0",x"c0",x"a0",x"80",x"60",x"ad",x"ff",x"ff",x"db",x"ff",x"d2",x"80",x"c0",x"c0",x"e0",x"e0",x"e0",x"c0",x"80",x"60",x"89",x"fb",x"ff",x"b6",x"00",x"00",x"00",x"00",x"00",x"00",x"92",x"fb",x"a9",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"80",x"88",x"d2",x"a0",x"c0",x"c0",x"a0",x"a0",x"80",x"64",x"92",x"ff",x"ff",x"b2",x"6e",x"ff",x"d6",x"84",x"a0",x"c0",x"c0",x"c0",x"c0",x"a0",x"80",x"60",x"b2",x"ff",x"ff",x"b7",x"25",x"bb",x"fb",x"a4",x"80",x"c0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"6d",x"db",x"ff",x"db",x"49",x"00",x"00",x"00",x"00",x"49",x"fb",x"ed",x"c0",x"e0",x"a0",x"64",x"ff",x"db",x"24",x"00",x"04",x"49",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"24",x"00",x"92",x"b2",x"60",x"80",x"80",x"80",x"80",x"80",x"a0",x"a4",x"f2",x"f6",x"ed",x"c4",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"e5",x"ed",x"f2",x"f6",x"f6",x"fb",x"fb",x"6e",x"6e",x"ff",x"db",x"89",x"80",x"80",x"60",x"64",x"8d",x"b6",x"ff",x"ff",x"d7",x"24",x"92",x"ff",x"b2",x"84",x"80",x"a0",x"a0",x"80",x"60",x"69",x"b2",x"ff",x"ff",x"b7",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"ff",x"d6",x"89",x"80",x"80",x"80",x"80",x"60",x"69",x"db",x"ff",x"a9",x"80",x"80",x"60",x"64",x"8d",x"db",x"ff",x"ff",x"b2",x"00",x"00",x"92",x"ff",x"d6",x"84",x"80",x"80",x"60",x"60",x"64",x"89",x"db",x"ff",x"ff",x"b6",x"20",x"00",x"4d",x"ff",x"fb",x"89",x"60",x"80",x"80",x"60",x"60",x"69",x"b6",x"ff",x"ff",x"bb",x"25",x"00",x"00",x"00",x"00",x"6a",x"f7",x"ee",x"c0",x"e0",x"c0",x"60",x"d6",x"ff",x"6e",x"00",x"00",x"24",x"6d",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"24",x"00",x"b7",x"d7",x"ad",x"b1",x"b2",x"b1",x"b2",x"b1",x"cd",x"ed",x"ed",x"e4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c4",x"c4",x"e9",x"ed",x"f6",x"fb",x"fb",x"ff",x"ff",x"fb",x"b2",x"b2",x"b2",x"db",x"ff",x"ff",x"ff",x"92",x"20",x"00",x"25",x"df",x"ff",x"f6",x"b1",x"8d",x"69",x"8d",x"b6",x"db",x"ff",x"ff",x"96",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"92",x"ff",x"fb",x"d2",x"ad",x"89",x"8d",x"b2",x"db",x"ff",x"ff",x"fb",x"b2",x"b2",x"b6",x"fb",x"ff",x"ff",x"df",x"92",x"00",x"00",x"00",x"25",x"db",x"ff",x"fb",x"d6",x"b2",x"b2",x"b6",x"db",x"ff",x"ff",x"ff",x"92",x"00",x"00",x"00",x"00",x"92",x"ff",x"ff",x"d6",x"b2",x"8d",x"b2",x"d6",x"ff",x"ff",x"ff",x"b6",x"25",x"00",x"00",x"00",x"00",x"69",x"f7",x"ee",x"c0",x"e0",x"c0",x"80",x"8d",x"ff",x"bb",x"00",x"00",x"04",x"49",x"92",x"92",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"49",x"00",x"00",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"f6",x"e9",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"c9",x"f2",x"f6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"d7",x"49",x"00",x"00",x"00",x"00",x"49",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"6e",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"b7",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"b7",x"b7",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"b7",x"25",x"00",x"00",x"00",x"00",x"00",x"29",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"bb",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"92",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"6e",x"00",x"00",x"00",x"00",x"00",x"6e",x"fb",x"ed",x"c0",x"e0",x"e0",x"a0",x"84",x"fb",x"ff",x"29",x"00",x"00",x"24",x"6d",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"49",x"00",x"05",x"db",x"ff",x"db",x"fb",x"ff",x"ff",x"fb",x"ee",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c4",x"e9",x"f2",x"fb",x"ff",x"ff",x"ff",x"92",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"29",x"b7",x"ff",x"ff",x"ff",x"ff",x"df",x"b7",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"6e",x"db",x"ff",x"ff",x"ff",x"ff",x"92",x"25",x"25",x"b7",x"ff",x"db",x"db",x"b7",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"92",x"db",x"ff",x"ff",x"db",x"b7",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6e",x"db",x"db",x"df",x"ff",x"b7",x"6e",x"25",x"00",x"00",x"00",x"00",x"25",x"b2",x"f7",x"ed",x"c0",x"e0",x"e0",x"c0",x"60",x"b6",x"ff",x"92",x"00",x"00",x"24",x"49",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"49",x"00",x"00",x"25",x"49",x"25",x"49",x"db",x"fb",x"e9",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c4",x"c9",x"f2",x"f6",x"fb",x"fb",x"b7",x"6e",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"49",x"6d",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"49",x"6d",x"6d",x"25",x"00",x"00",x"00",x"00",x"25",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"25",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"05",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"d7",x"f7",x"c9",x"c0",x"e0",x"e0",x"c0",x"60",x"b2",x"ff",x"d7",x"24",x"00",x"24",x"49",x"6d",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"6d",x"29",x"00",x"00",x"00",x"00",x"00",x"92",x"fb",x"e9",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e9",x"f2",x"f6",x"fb",x"fb",x"b6",x"6e",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"b2",x"fb",x"f2",x"c4",x"c0",x"e0",x"e0",x"c0",x"60",x"8d",x"ff",x"db",x"49",x"00",x"00",x"24",x"49",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"6d",x"29",x"00",x"00",x"00",x"00",x"6e",x"fb",x"c9",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c4",x"cd",x"f2",x"fb",x"fb",x"fb",x"b6",x"6e",x"29",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"fb",x"f7",x"e9",x"c0",x"e0",x"e0",x"e0",x"c0",x"60",x"89",x"db",x"df",x"4d",x"00",x"00",x"24",x"49",x"6d",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"92",x"6d",x"25",x"00",x"00",x"00",x"6e",x"fb",x"cd",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c4",x"c9",x"d2",x"f7",x"fb",x"db",x"b7",x"b2",x"69",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"6e",x"d7",x"f7",x"f2",x"c5",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"69",x"db",x"ff",x"72",x"00",x"00",x"24",x"24",x"6d",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"49",x"24",x"00",x"00",x"25",x"fb",x"f2",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a4",x"a9",x"cd",x"d2",x"f7",x"d7",x"d7",x"b6",x"92",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"92",x"d7",x"f7",x"f2",x"e9",x"c0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"64",x"db",x"ff",x"b6",x"00",x"00",x"00",x"49",x"6d",x"6d",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"49",x"00",x"00",x"00",x"d7",x"f2",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"84",x"84",x"88",x"ad",x"b2",x"b2",x"b2",x"b2",x"8e",x"69",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"6d",x"b2",x"d7",x"f7",x"f2",x"c5",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"89",x"d7",x"ff",x"b7",x"24",x"00",x"00",x"24",x"49",x"6d",x"b6",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"6d",x"24",x"00",x"00",x"6e",x"fb",x"c5",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"64",x"69",x"89",x"8e",x"b2",x"92",x"92",x"6e",x"6e",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"6d",x"92",x"db",x"fb",x"f7",x"f2",x"e9",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"60",x"68",x"da",x"ff",x"db",x"25",x"00",x"00",x"24",x"49",x"6d",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"6e",x"49",x"24",x"00",x"49",x"db",x"e9",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"64",x"64",x"45",x"69",x"8d",x"8e",x"8e",x"6e",x"6d",x"4d",x"49",x"49",x"25",x"25",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"69",x"6e",x"92",x"b7",x"d7",x"d7",x"f6",x"f2",x"ed",x"c5",x"e0",x"e0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"60",x"89",x"db",x"ff",x"b7",x"45",x"00",x"00",x"24",x"49",x"6d",x"92",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"6d",x"24",x"00",x"00",x"b2",x"f7",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"60",x"40",x"40",x"40",x"40",x"64",x"65",x"69",x"69",x"8d",x"8d",x"8e",x"8e",x"6e",x"6e",x"6e",x"6d",x"49",x"49",x"49",x"49",x"29",x"29",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"29",x"49",x"49",x"49",x"6e",x"92",x"92",x"b6",x"d7",x"f7",x"fb",x"fb",x"f7",x"f2",x"e9",x"c5",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"60",x"8d",x"db",x"ff",x"b7",x"25",x"00",x"00",x"24",x"49",x"6d",x"92",x"b6",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"49",x"24",x"00",x"49",x"f7",x"c5",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"40",x"60",x"60",x"80",x"80",x"80",x"80",x"a4",x"a4",x"a4",x"a4",x"a4",x"c4",x"c4",x"a8",x"a4",x"c4",x"a4",x"a4",x"a4",x"a4",x"a4",x"84",x"84",x"80",x"80",x"60",x"64",x"64",x"64",x"65",x"69",x"69",x"89",x"8d",x"92",x"92",x"92",x"b2",x"b2",x"b2",x"b2",x"b2",x"b2",x"b2",x"b6",x"b6",x"b6",x"b7",x"b7",x"b7",x"b7",x"b7",x"d7",x"d7",x"fb",x"f7",x"f7",x"fb",x"f7",x"f6",x"f2",x"ee",x"ed",x"e9",x"e5",x"c0",x"e0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"64",x"b1",x"ff",x"ff",x"b7",x"25",x"00",x"00",x"20",x"24",x"49",x"6d",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"92",x"6d",x"45",x"00",x"00",x"b7",x"f2",x"e0",x"e0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"60",x"60",x"60",x"80",x"84",x"a4",x"c4",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c8",x"e8",x"e8",x"ec",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"c4",x"a4",x"84",x"60",x"60",x"60",x"40",x"40",x"44",x"64",x"69",x"89",x"a9",x"ad",x"ae",x"ce",x"d2",x"f6",x"f6",x"f6",x"f6",x"f6",x"f7",x"f7",x"f6",x"f2",x"f2",x"f2",x"ee",x"ee",x"ed",x"e9",x"e5",x"e5",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"80",x"64",x"b6",x"ff",x"ff",x"b6",x"25",x"00",x"00",x"24",x"24",x"49",x"6d",x"92",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"49",x"24",x"00",x"49",x"fb",x"c5",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"80",x"60",x"60",x"60",x"40",x"60",x"60",x"80",x"a4",x"a4",x"c4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c8",x"c8",x"e8",x"e8",x"e8",x"e8",x"e4",x"cc",x"cc",x"e8",x"e8",x"e8",x"e8",x"e8",x"c8",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"c4",x"a0",x"80",x"60",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"80",x"a0",x"a4",x"c4",x"c4",x"c4",x"c4",x"c4",x"c4",x"c0",x"e0",x"c0",x"c0",x"e0",x"e0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"60",x"89",x"db",x"ff",x"df",x"92",x"00",x"00",x"00",x"24",x"48",x"49",x"6d",x"92",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"6e",x"49",x"00",x"00",x"b2",x"f2",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"80",x"a4",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e4",x"e4",x"c8",x"c8",x"e4",x"e4",x"e8",x"c4",x"cc",x"f6",x"fa",x"f6",x"e8",x"e4",x"c8",x"d1",x"d6",x"f6",x"ec",x"e4",x"e8",x"c8",x"c8",x"e8",x"e8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"c4",x"a4",x"80",x"60",x"60",x"40",x"60",x"60",x"80",x"a0",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"64",x"b1",x"ff",x"ff",x"db",x"6e",x"00",x"00",x"00",x"24",x"48",x"49",x"6d",x"92",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"24",x"00",x"25",x"f7",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a0",x"80",x"80",x"64",x"89",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"89",x"69",x"88",x"84",x"84",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"60",x"60",x"60",x"a0",x"c4",x"c8",x"e8",x"e8",x"e8",x"e8",x"c8",x"e8",x"e4",x"e4",x"e4",x"e4",x"e4",x"c8",x"f6",x"f6",x"e8",x"e4",x"e4",x"c8",x"f6",x"ff",x"ff",x"ff",x"f1",x"e4",x"cd",x"ff",x"ff",x"ff",x"f6",x"e4",x"e8",x"f1",x"f1",x"e4",x"e4",x"e4",x"c8",x"c8",x"c8",x"c8",x"e8",x"e8",x"e8",x"e8",x"c4",x"a4",x"80",x"60",x"60",x"60",x"80",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"60",x"8d",x"db",x"ff",x"ff",x"b7",x"49",x"00",x"00",x"00",x"24",x"48",x"49",x"6d",x"92",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"49",x"24",x"00",x"6e",x"f2",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"69",x"b2",x"d6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"db",x"d6",x"d6",x"ae",x"89",x"64",x"60",x"80",x"80",x"80",x"a0",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"80",x"a0",x"c4",x"e8",x"e8",x"e8",x"e4",x"e4",x"e4",x"c8",x"ac",x"c8",x"e4",x"e4",x"e4",x"e4",x"e4",x"cd",x"ff",x"ff",x"ed",x"e4",x"e4",x"c9",x"ff",x"ff",x"f6",x"ff",x"f1",x"e4",x"f2",x"ff",x"fb",x"ff",x"fa",x"e4",x"e8",x"ff",x"f6",x"e4",x"c4",x"c8",x"d1",x"f6",x"f6",x"d1",x"c8",x"e4",x"e4",x"e8",x"e8",x"e8",x"e8",x"a4",x"80",x"80",x"80",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"60",x"64",x"b6",x"ff",x"ff",x"ff",x"92",x"00",x"00",x"00",x"00",x"24",x"49",x"6d",x"6d",x"92",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"6d",x"49",x"20",x"00",x"d7",x"c9",x"e0",x"e0",x"e0",x"e0",x"a0",x"80",x"84",x"8d",x"db",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"b2",x"ad",x"89",x"84",x"80",x"a0",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"a0",x"c8",x"e8",x"e8",x"e4",x"c4",x"cd",x"f1",x"f1",x"c4",x"c9",x"ff",x"f1",x"e0",x"e4",x"e4",x"e4",x"e4",x"f2",x"ff",x"ff",x"f2",x"c4",x"e0",x"c9",x"ff",x"f6",x"e5",x"ed",x"c8",x"c4",x"f7",x"ff",x"cd",x"d1",x"f2",x"e4",x"e8",x"ff",x"f6",x"e4",x"c4",x"d1",x"ff",x"ff",x"ff",x"fb",x"ed",x"e4",x"e4",x"c8",x"c8",x"c8",x"e8",x"e8",x"e8",x"a4",x"80",x"80",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"64",x"b6",x"df",x"ff",x"ff",x"b7",x"49",x"00",x"00",x"00",x"04",x"24",x"49",x"6d",x"6e",x"92",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"24",x"00",x"49",x"f7",x"e4",x"e0",x"e0",x"c0",x"80",x"40",x"6d",x"db",x"ff",x"ff",x"ff",x"ff",x"db",x"b7",x"92",x"6e",x"4d",x"49",x"49",x"49",x"49",x"6e",x"6e",x"92",x"b6",x"b7",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"db",x"d6",x"ae",x"89",x"60",x"60",x"80",x"80",x"c0",x"c0",x"e0",x"e0",x"c0",x"a0",x"60",x"c4",x"e4",x"e4",x"e4",x"c4",x"d1",x"fb",x"ff",x"ff",x"cd",x"ed",x"ff",x"ed",x"e0",x"e4",x"e4",x"e4",x"e0",x"f6",x"ff",x"ff",x"f7",x"c4",x"e0",x"cd",x"ff",x"d1",x"a0",x"e4",x"c4",x"c4",x"fb",x"ff",x"c8",x"e0",x"e4",x"e4",x"e4",x"ff",x"fa",x"e4",x"e4",x"fb",x"ff",x"fb",x"ff",x"ff",x"fa",x"c4",x"c8",x"d6",x"fb",x"f2",x"c4",x"e4",x"e4",x"e4",x"60",x"80",x"a0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"80",x"60",x"68",x"b6",x"db",x"ff",x"ff",x"db",x"8e",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"6d",x"92",x"92",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"b6",x"92",x"49",x"24",x"00",x"92",x"ee",x"e0",x"e0",x"c0",x"80",x"64",x"d6",x"ff",x"ff",x"ff",x"db",x"6e",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"8e",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"b2",x"8d",x"68",x"64",x"60",x"80",x"80",x"60",x"40",x"a4",x"e4",x"e4",x"c4",x"cc",x"ff",x"ff",x"ff",x"ff",x"ed",x"ed",x"ff",x"ed",x"e0",x"e4",x"e4",x"e4",x"e4",x"fb",x"fb",x"fb",x"ff",x"c4",x"e0",x"ed",x"ff",x"fb",x"cd",x"c4",x"e0",x"e0",x"f6",x"ff",x"f2",x"c4",x"e0",x"e0",x"e8",x"ff",x"f6",x"c4",x"c9",x"ff",x"fb",x"ed",x"cd",x"fa",x"f6",x"c4",x"f2",x"ff",x"ff",x"ff",x"f2",x"e4",x"e4",x"e4",x"60",x"80",x"a0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"80",x"60",x"60",x"8d",x"d6",x"fb",x"ff",x"ff",x"db",x"6e",x"24",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"6d",x"92",x"92",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"49",x"00",x"00",x"d6",x"e9",x"e0",x"c0",x"60",x"89",x"db",x"ff",x"ff",x"bb",x"6e",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"6d",x"92",x"b7",x"db",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"b2",x"89",x"64",x"20",x"20",x"a4",x"e4",x"e0",x"c4",x"d6",x"ff",x"fb",x"f6",x"fa",x"e8",x"ed",x"ff",x"ed",x"e0",x"e4",x"e4",x"e0",x"c8",x"ff",x"d2",x"f6",x"ff",x"ed",x"e0",x"c8",x"fb",x"ff",x"fb",x"cd",x"e0",x"e0",x"f2",x"ff",x"ff",x"d2",x"c4",x"e0",x"e8",x"ff",x"f6",x"c4",x"f1",x"ff",x"f2",x"c0",x"c4",x"e9",x"ed",x"c4",x"f6",x"ff",x"fb",x"ff",x"fb",x"e0",x"e4",x"e4",x"80",x"80",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"40",x"40",x"8d",x"b6",x"df",x"ff",x"ff",x"fb",x"b2",x"49",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"6d",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"6d",x"24",x"00",x"25",x"f7",x"c0",x"a0",x"60",x"b2",x"ff",x"ff",x"db",x"4d",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"04",x"24",x"24",x"24",x"04",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"92",x"b7",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"d7",x"8e",x"49",x"a4",x"e4",x"e0",x"c9",x"ff",x"fa",x"c4",x"c0",x"c4",x"e0",x"ed",x"ff",x"ed",x"e0",x"e4",x"e4",x"e0",x"cd",x"ff",x"cd",x"ed",x"ff",x"ed",x"e0",x"e0",x"ed",x"ff",x"ff",x"fb",x"ed",x"e0",x"c4",x"f6",x"ff",x"ff",x"f2",x"c0",x"e4",x"ff",x"fa",x"e0",x"f2",x"ff",x"cd",x"c0",x"e0",x"e0",x"e0",x"c0",x"fb",x"ff",x"a5",x"cd",x"f6",x"e0",x"e4",x"e4",x"60",x"60",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"60",x"84",x"ad",x"d6",x"fb",x"ff",x"ff",x"ff",x"db",x"6e",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"6d",x"6d",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"24",x"00",x"8e",x"f2",x"a0",x"60",x"b2",x"ff",x"ff",x"b7",x"25",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"48",x"48",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"29",x"6d",x"92",x"b7",x"df",x"ff",x"ff",x"bb",x"92",x"a4",x"e0",x"e0",x"cd",x"ff",x"ed",x"e0",x"e0",x"e0",x"e0",x"ed",x"ff",x"ed",x"e0",x"e0",x"e4",x"e0",x"f2",x"ff",x"a5",x"c9",x"ff",x"f2",x"e0",x"e0",x"e4",x"cd",x"fb",x"ff",x"f6",x"c0",x"e0",x"c8",x"f6",x"ff",x"ff",x"c4",x"e4",x"ff",x"fa",x"c0",x"f2",x"ff",x"cd",x"e0",x"e0",x"e0",x"e0",x"e0",x"f6",x"ff",x"c9",x"c0",x"e4",x"e0",x"e4",x"e4",x"60",x"60",x"a0",x"c0",x"c0",x"e0",x"e0",x"c0",x"a0",x"a0",x"80",x"60",x"40",x"64",x"b1",x"d6",x"fb",x"ff",x"ff",x"ff",x"ff",x"db",x"8e",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"49",x"00",x"00",x"d7",x"a9",x"60",x"b2",x"ff",x"ff",x"6e",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"4d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"25",x"49",x"4d",x"6d",x"a4",x"e0",x"e0",x"f6",x"ff",x"c8",x"e0",x"e0",x"e0",x"e0",x"ed",x"ff",x"ed",x"e0",x"e0",x"e0",x"c0",x"fa",x"ff",x"b1",x"d2",x"ff",x"fb",x"c4",x"e0",x"e0",x"c0",x"e9",x"ff",x"fa",x"e0",x"e0",x"e0",x"c4",x"f7",x"ff",x"e9",x"e4",x"ff",x"f6",x"c0",x"f2",x"ff",x"c9",x"e0",x"e0",x"e0",x"e0",x"e0",x"ed",x"ff",x"f6",x"c0",x"e0",x"e0",x"e0",x"e0",x"40",x"40",x"80",x"80",x"80",x"80",x"60",x"60",x"64",x"89",x"ad",x"d2",x"d6",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"29",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"48",x"49",x"49",x"6d",x"6d",x"92",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"b6",x"92",x"49",x"00",x"24",x"d7",x"64",x"8d",x"ff",x"ff",x"6e",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"91",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"e0",x"e4",x"fb",x"fb",x"c4",x"e0",x"e0",x"e0",x"e0",x"ed",x"ff",x"ed",x"e0",x"e0",x"e0",x"c4",x"ff",x"ff",x"fb",x"ff",x"ff",x"fb",x"c9",x"c0",x"c0",x"c0",x"c4",x"ff",x"fb",x"e0",x"c0",x"e4",x"a0",x"d2",x"ff",x"ed",x"e4",x"ff",x"f6",x"c0",x"f2",x"ff",x"ed",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"fa",x"ff",x"f2",x"c0",x"e0",x"e0",x"c0",x"20",x"20",x"20",x"60",x"64",x"89",x"ad",x"b2",x"d6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"96",x"6d",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"49",x"00",x"49",x"b2",x"69",x"db",x"ff",x"6e",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"e0",x"e4",x"fb",x"fb",x"e0",x"e0",x"e0",x"e0",x"e0",x"ed",x"ff",x"ed",x"e0",x"e0",x"e0",x"c9",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"c9",x"c4",x"f2",x"e9",x"cd",x"ff",x"f7",x"c0",x"ed",x"f1",x"a4",x"d6",x"ff",x"cd",x"c4",x"ff",x"f7",x"e0",x"ed",x"ff",x"f2",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"ed",x"ff",x"ff",x"ed",x"e0",x"e0",x"c0",x"44",x"49",x"6e",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"bb",x"92",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"24",x"00",x"92",x"b6",x"db",x"ff",x"92",x"00",x"00",x"00",x"00",x"24",x"49",x"6d",x"6d",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"8e",x"6d",x"6d",x"6d",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"e0",x"c4",x"fb",x"fb",x"c4",x"e0",x"e0",x"c0",x"e0",x"ed",x"ff",x"cd",x"a4",x"e4",x"c0",x"cd",x"ff",x"d6",x"cd",x"c9",x"d6",x"ff",x"cd",x"c9",x"ff",x"fb",x"fb",x"ff",x"ee",x"c0",x"f6",x"ff",x"f7",x"ff",x"ff",x"c4",x"c4",x"ff",x"f6",x"e0",x"c4",x"ff",x"fb",x"c8",x"c0",x"c0",x"c0",x"e0",x"e0",x"c0",x"ee",x"ff",x"fb",x"c4",x"e0",x"c0",x"69",x"72",x"97",x"bb",x"db",x"df",x"db",x"b7",x"b2",x"92",x"49",x"45",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"d7",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"48",x"00",x"92",x"ff",x"ff",x"b7",x"00",x"00",x"00",x"00",x"24",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"80",x"e0",x"e0",x"fb",x"ff",x"c4",x"e0",x"c0",x"e4",x"e0",x"ed",x"ff",x"f6",x"f2",x"f6",x"c4",x"f2",x"ff",x"c9",x"e0",x"c0",x"c9",x"ff",x"d1",x"c9",x"ff",x"ff",x"ff",x"fb",x"e9",x"c0",x"f6",x"ff",x"ff",x"ff",x"fb",x"c0",x"c4",x"ff",x"f6",x"e0",x"c0",x"f6",x"ff",x"f6",x"c9",x"cd",x"ed",x"e0",x"c0",x"c0",x"c0",x"f6",x"ff",x"e9",x"e0",x"c0",x"64",x"4d",x"4d",x"49",x"49",x"49",x"25",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"49",x"00",x"25",x"db",x"db",x"25",x"00",x"00",x"00",x"24",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"6d",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"a0",x"e0",x"e0",x"fb",x"ff",x"ed",x"c0",x"c9",x"f6",x"e9",x"cd",x"ff",x"ff",x"ff",x"ff",x"e9",x"f6",x"fb",x"e4",x"e0",x"e0",x"e4",x"f2",x"e9",x"c4",x"ee",x"f6",x"f2",x"e9",x"e0",x"e0",x"e9",x"f6",x"fb",x"f6",x"e9",x"e0",x"e0",x"f6",x"f2",x"c0",x"e0",x"ed",x"ff",x"ff",x"fb",x"ff",x"f6",x"c0",x"c9",x"c9",x"a0",x"ce",x"ff",x"e9",x"e0",x"c0",x"40",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"b6",x"92",x"49",x"00",x"00",x"49",x"49",x"00",x"00",x"00",x"24",x"49",x"6d",x"92",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"92",x"69",x"24",x"00",x"00",x"00",x"20",x"40",x"40",x"40",x"a0",x"e0",x"e0",x"f2",x"ff",x"fb",x"d2",x"da",x"ff",x"cd",x"cd",x"ff",x"ff",x"fb",x"f6",x"e4",x"ed",x"ed",x"e0",x"e0",x"e0",x"e0",x"e4",x"e0",x"e0",x"e0",x"c4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e4",x"c9",x"c4",x"e0",x"e0",x"e0",x"e5",x"e4",x"c0",x"e0",x"e0",x"f2",x"ff",x"ff",x"ff",x"f6",x"c0",x"f6",x"f6",x"c9",x"d6",x"ff",x"ed",x"e0",x"c0",x"40",x"40",x"40",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"6d",x"92",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"92",x"6d",x"24",x"00",x"20",x"40",x"80",x"a0",x"80",x"40",x"a0",x"e0",x"e0",x"cd",x"ff",x"ff",x"ff",x"ff",x"fb",x"c8",x"e8",x"f2",x"cd",x"cd",x"c4",x"e0",x"e0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"e0",x"e0",x"e0",x"c4",x"f2",x"fb",x"f6",x"e9",x"c0",x"f6",x"ff",x"fb",x"ff",x"ff",x"e9",x"e0",x"c0",x"60",x"60",x"a0",x"80",x"40",x"20",x"00",x"00",x"24",x"24",x"29",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"6d",x"49",x"00",x"00",x"00",x"00",x"24",x"49",x"6d",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"96",x"6d",x"24",x"00",x"60",x"a0",x"c0",x"e0",x"a0",x"60",x"a0",x"e0",x"e0",x"c4",x"f6",x"ff",x"ff",x"fb",x"ee",x"c0",x"e0",x"e0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"e0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"c5",x"e0",x"e0",x"e9",x"fb",x"ff",x"ff",x"fb",x"e4",x"e0",x"c0",x"60",x"80",x"a0",x"c0",x"c0",x"80",x"20",x"00",x"24",x"49",x"49",x"6d",x"6d",x"91",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"6d",x"49",x"24",x"24",x"48",x"49",x"6d",x"92",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"72",x"45",x"20",x"a4",x"e0",x"e0",x"c0",x"80",x"60",x"a0",x"e0",x"e0",x"e0",x"e5",x"ee",x"f2",x"e9",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"e0",x"e0",x"e0",x"ed",x"f6",x"f7",x"ed",x"c0",x"e0",x"c0",x"60",x"80",x"a0",x"e0",x"e0",x"c0",x"40",x"00",x"24",x"49",x"6d",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"6d",x"49",x"49",x"6d",x"6d",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"49",x"00",x"80",x"e0",x"e0",x"c0",x"80",x"60",x"a0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"80",x"80",x"40",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"40",x"60",x"80",x"80",x"a0",x"c0",x"c0",x"e0",x"e4",x"e0",x"e0",x"c0",x"c0",x"e5",x"c0",x"e0",x"e0",x"e0",x"60",x"80",x"c0",x"e0",x"e0",x"c0",x"40",x"00",x"48",x"6d",x"92",x"b6",x"b6",x"b7",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"92",x"71",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"49",x"00",x"40",x"c0",x"e0",x"c0",x"80",x"40",x"a0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a4",x"a4",x"60",x"60",x"40",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"40",x"60",x"60",x"a0",x"a4",x"c0",x"e0",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"40",x"60",x"c0",x"e0",x"e0",x"80",x"20",x"24",x"49",x"6d",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"b6",x"92",x"92",x"92",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"49",x"20",x"00",x"60",x"e0",x"c0",x"80",x"40",x"a0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"84",x"60",x"40",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"60",x"84",x"a4",x"c0",x"e0",x"e0",x"e0",x"e0",x"c0",x"60",x"60",x"a0",x"e0",x"a0",x"20",x"00",x"24",x"6d",x"92",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"49",x"24",x"00",x"20",x"a0",x"c0",x"a0",x"60",x"a0",x"c0",x"c0",x"c4",x"a0",x"60",x"40",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"40",x"60",x"80",x"a0",x"c0",x"e0",x"c0",x"60",x"80",x"a0",x"c0",x"60",x"00",x"00",x"24",x"6d",x"92",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"49",x"24",x"00",x"00",x"60",x"c0",x"a0",x"60",x"84",x"a4",x"80",x"40",x"20",x"00",x"00",x"00",x"00",x"04",x"24",x"24",x"24",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"04",x"04",x"00",x"00",x"00",x"00",x"20",x"40",x"80",x"a0",x"a4",x"60",x"80",x"a0",x"a0",x"20",x"00",x"00",x"49",x"6d",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"24",x"00",x"00",x"60",x"c0",x"a0",x"40",x"40",x"40",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"28",x"29",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"24",x"04",x"04",x"00",x"00",x"00",x"00",x"20",x"40",x"40",x"60",x"c0",x"a0",x"00",x"00",x"20",x"49",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"24",x"00",x"00",x"60",x"c0",x"80",x"40",x"00",x"00",x"00",x"00",x"20",x"24",x"44",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"69",x"69",x"49",x"49",x"29",x"24",x"04",x"00",x"00",x"00",x"20",x"20",x"60",x"c0",x"a0",x"00",x"00",x"24",x"49",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"24",x"00",x"20",x"a0",x"c0",x"80",x"40",x"00",x"00",x"00",x"20",x"24",x"49",x"49",x"6d",x"6d",x"8d",x"8e",x"92",x"92",x"96",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"72",x"6d",x"6d",x"6d",x"49",x"49",x"24",x"24",x"00",x"00",x"20",x"40",x"80",x"c0",x"c0",x"40",x"00",x"24",x"49",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"24",x"00",x"40",x"c0",x"e0",x"80",x"40",x"00",x"00",x"00",x"44",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"b2",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"96",x"92",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"24",x"00",x"00",x"20",x"80",x"c0",x"e0",x"60",x"00",x"00",x"49",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"24",x"00",x"80",x"e0",x"e0",x"80",x"60",x"20",x"00",x"24",x"49",x"6d",x"92",x"92",x"b2",x"b6",x"b6",x"b7",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"d7",x"b6",x"b6",x"96",x"92",x"92",x"6d",x"49",x"24",x"04",x"00",x"20",x"60",x"a0",x"e0",x"a0",x"00",x"00",x"49",x"6d",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"69",x"00",x"20",x"a0",x"e0",x"e0",x"a0",x"40",x"00",x"24",x"49",x"6d",x"92",x"b2",x"b6",x"b6",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"6d",x"49",x"24",x"00",x"20",x"60",x"c0",x"e0",x"c0",x"20",x"00",x"28",x"6d",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"49",x"00",x"40",x"c0",x"e0",x"c0",x"60",x"20",x"00",x"24",x"49",x"92",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"92",x"6d",x"49",x"00",x"00",x"40",x"c0",x"e0",x"e0",x"80",x"00",x"24",x"8d",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"db",x"92",x"49",x"00",x"80",x"c0",x"a0",x"60",x"20",x"00",x"24",x"49",x"6d",x"92",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"6d",x"49",x"24",x"00",x"20",x"60",x"c0",x"c0",x"a0",x"20",x"24",x"6d",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"d6",x"92",x"49",x"00",x"80",x"80",x"40",x"20",x"00",x"04",x"44",x"6d",x"92",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"6d",x"49",x"20",x"00",x"00",x"40",x"80",x"a4",x"40",x"24",x"6d",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"49",x"00",x"40",x"20",x"00",x"00",x"24",x"45",x"49",x"92",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"92",x"4d",x"48",x"24",x"00",x"00",x"20",x"40",x"20",x"24",x"71",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"96",x"6d",x"20",x"00",x"00",x"00",x"04",x"49",x"49",x"6d",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"92",x"6d",x"4d",x"48",x"24",x"00",x"00",x"00",x"00",x"24",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"8d",x"49",x"24",x"24",x"24",x"49",x"4d",x"6d",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"6d",x"6d",x"49",x"24",x"24",x"00",x"20",x"49",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"92",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"8e",x"6d",x"49",x"49",x"49",x"49",x"6d",x"b6",x"db",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"db",x"96",x"92",x"6d",x"6d",x"6d",x"92",x"92",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"92",x"72",x"6d",x"6d",x"6d",x"6d",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"b6",x"92",x"92",x"92",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"92",x"92",x"92",x"92",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff")
);
	constant logo1_Mask : mask_array := (
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111100000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000001111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111100000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000011111111111111111111111110000000000000000000000000000000111110000000000000000000000000000000000000011111111111101111110000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000011111111111111111111111111111111111111000000000000000001111111000000000000000000111111111111100000111111111111101111111000000000001111111000000000111111110000000000000000000000000000"),
("00000000000000000011111111111111111111111111111111111111111000000000000011111111000000000000000001111111111111110001111111111111001111111100000001111111111111000011111111111000000000000000000000000000"),
("00000000000000000011111111111111111111111111111111111111111100000000000111111111110000000000000011111111111111111101111111111111001111111110000011111111111111111111111111111110000000000000000000000000"),
("00000000000000000011111011111111111111111111111111111111111111000000000111111111110000000000000111111111111111111111111111111111001111111111111111111111111111111111111111111111000000000000000000000000"),
("00000000000000000011111011111111111111111111111111111111111111100000001111111111111000000000000111111111111111111111111111111110000111111111111111111111111111111111111111111111000000000000000000000000"),
("00000000000000000011111011111111111111111111111111111111111111100000011111111111111100000000000111111111111111111111111111111110000111111111111111111111111111111111111111111111100000000000000000000000"),
("00000000000000000011111111111111111111111111111111111111111111110000111111111111111110000000001111111111111111111111111111011100000111111111111111111111111111111111111111111111110000000000000000000000"),
("00000000000000000011111111111111111111111111111111111111111111111000111111111111111111000000001111111111111111111111111110000000000111111111111111111111111111111111111111111111110000000000000000000000"),
("00000000000000000011111111111111111111111111111111111111111111111111111111110111111111000000001111111111111111111111111111000000000011111111111111111111111111111111111111111111110000000000000000000000"),
("00000000000000000011111101111111111111110011111111111111111111111111111111110111111111100000001111111111111111111111111111000000000000011111111111111111111111111111111111111111111000000000000000000000"),
("00000000000000000011111111111111111111111111111111111111111111111111111111100111111111100000011111110111111101111111111111100000000000000111111111111111111111111111111111111111111000000000000000000000"),
("00000000000000000011111110111111111111111111111111111111111111111111111111100111111111100000011111101111111111111111111111110000000000001111111111111111111111111110111111111111111000000000000000000000"),
("00000000000000000111111110111111111111111111111111111111111111111111111100000000111111110000011111111111111111111111111111110000000000001111111111111111111111111111111111111111111000000000000000000000"),
("00000000000000011111111111011111111111111111111111111111111111111111111100000000111111110000111111111111111101111111111111111000000000011111111111111111111111111011111111111111111100000000000000000000"),
("00000000000000111111111111101111111111111111111111111111111111111111111110000001111111111000111111111111111111111111111111111000000000111111111111111111111111110111111111111111111100000000000000000000"),
("00000000000001111111111111110001111111111111111111111111111111111111111110000001111111111000111111011111111111111111111111111000000001111111111011111111111111111111111111111111111100000000000000000000"),
("00000000000011111111111111111100011111111111111111111111111111111111111111000011111111111000111111111111111111111111111111110000000001111111111111111111111111011111111111111111111100000000000000000000"),
("00000000000011111111111111111111100111111111111101111111111111111111111111000011111111111101111111111111111011111111111111110000000001111111110111111111111111011111111111111111111100000000000000000000"),
("00000000000111111111111111111111111011111111111000011111111111111111111110000011111111111111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111100000000000000000000"),
("00000000000111111111111111111111111111111111110111111111111101111111111110010011111111111111111111111111111111111111111111110000000001111111101111111110111110111111111011111111111100000000000000000000"),
("00000000001111111111111111111111111111111111110111111111111101110111111110111011111111111111111111111111111111111111111111110001100001111111111111111110111110111111111011111111111100000111100000000000"),
("00000000011111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111110111111111111111110011110001111111111111111101111111111111111011111011111100111111110000000000"),
("00000000111111111111111111111111111111111111111111011111111111011111111111111111111111111111111111111111111111111111111111100111111001111111111111111101111111111111110111111111111111111111111000000000"),
("00000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111101111111011111111101111101111111110111111111111111111111111100000000"),
("00000111111111101111111111111111111111111111111111111111111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111110111110111111111111111111110000000"),
("00000111111111101111111111111111111111111111011111111111111001111111111111111111111111111111111111111111101111111111111111111111111111111111111111111011111111111111110111110111111111111111111110000000"),
("00001111111111101111111111111111111111111111011111111111111011111111110111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111101111111111111111111111111111000000"),
("00001111111111000111111111111111111111111111111111111111111011111111111111111111111111111111111011111111111111111111111111111111111111111110111111111011111011111111101111111111111111111111111111100000"),
("00011111111111000111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111011111111101111101111111111111111111111110000"),
("00011111111110000111111111111111111111111111111111111111111111111111101111111111111111111111111111111111011111111111111111111111111111111111111111110111111111111111101111101111111111111111111111110000"),
("00011111111110000111111111111111111111111111111111111111111101111111011111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111011111111111111111111111111111110000"),
("00011111000000000000001111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111101111111110111110111111111011111111111111111111111111111111000"),
("00011111000000000000011111111111111111111111111111111111101110001001111111111111111111111111111111111110111111111111111111111111111111111111111111111111110111111111011111111111111111111111011111111000"),
("00011111100000000000011111111111111111111111111111111111111111100111111111111111111111111111111111111110111111111111111111111111111111111111111111101111111111111111111111111111111111111111011111111000"),
("00011111100000000000111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111110111111111111111111111100000011111000"),
("00011111110000000001111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111011111111101111111111111110111111111111111111111000000011111000"),
("00011111110000000011111111111111111111111111111111111111010111111111110111111111111111111111111111111101111111111111111111111111111111111111111111111111101111111110111111111111111111111100000111111000"),
("00011111111000000011111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111011111111111111111111111111111111111111100000111111000"),
("00001111111000000011111111111111111111111011111111111111111111111111111111111101111111111111111111111100011111111111111100001111111111111111111111011111011111111101111111111111111111111110000111111000"),
("00001111110000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111011111111111111101111111111111111110000111111000"),
("00001111110000000011111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111110000111111000"),
("00001111110000000011111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111101111111111111111110111111111111111011111111111111111110111011111000"),
("00001111110001100011111111111111111111110111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111101111111111111111110111111111111111011111111111111111110111111111000"),
("00011111110011100011111111111111111111111111111111111111111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111000"),
("00011111100111110011111111111111111111111111111111111101111111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111110111111111111111111111111111111000"),
("00011111101111111011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111111111001111111111111101111111111111111111111111111111000"),
("00011111111111111111111111111111111111101111111111111111111111111111111111111001111111111111111111110111111111111111111110111111111011111111111111110111111111111111101111111111111111111111111111111000"),
("00001111111111111111111111111111111111111111111111111011111111111111111111111011111111111111111111110111111111111111111110111111111111111111111111111111111111111111011111111111111111111111111111110000"),
("00001111111111111111111111111111111111111111111111111111111111110111111111111011111111111111111111110111111111111111111100111111111111111111111111101111111111111110111111111111111111111111111111110000"),
("00001111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111101111111111111111111101111111110111111111111111011111111111111100111111111111111111111111111111110000"),
("00001111111111111111111111111111111111011111111111110111111111111111111111110111111111111111111111101111111111111111111101111111110111111111111110111111111111111001111111111111111111111111111111100000"),
("00001111111111111111111111111111111111111111111111110111111111101111111111110111111111111111111111101111111111111111111101111111111111111111111101111111111111110011111111111111111111111111111111100000"),
("00001111111111111111111111111111111111111111111111101111111111111111111111110111111111111111111111101111111111111111111001111111111111111111111011111111111111100111111111111111111111111111111111000000"),
("00000111111111111111111111111111111111111111111111101111111111111111111111100111111111111111111111011111111111111111111011111111101111111111110111111111111111111111111111111100011111111111111100000000"),
("00000111111111111111111111111111111110111111111111011111111111111111111111101111111110111111111111011111111111111111111111111111111111111111111111111111111111011111111111111001111111111111111000000000"),
("00000011111111111111111111111111111110111111111111111111111111011111111111101111111110111111111111011111111011111111111111111111111111111111111111111111111111111111111111110111111111111111100000000000"),
("00000001111111111111111111111111111110111111111110111111111111011111111111101111111111111111111110011111111111111111110011111111111111111111111111111111111111111111111111101111111111111111000000000000"),
("00000000111111111111111111111111111111111111111101111111111111111111111111001111111111111111111110111111111111111111110111111111011111111111101111111111111111111111111111101111111111111110000000000000"),
("00000000001111111111111111111111111111111111111011111111111111111111111111011111111111111111111110111111110111111111110111111111011111111111111111111111111110111111111111011111111111111110000000000000"),
("00000000000001111111111111111111111111111111110111111111111110111111111111011111111111111111111110111111110111111111110111111111111111111111111111111111111111111111111111111111111111111110000000000000"),
("00000000000000011111111111111111111111111111100111111111111110111111111111011111111111111111111101111111111111111111100111111111111111111111011111111111111111111111111110111111111101111110000000000000"),
("00000000000000000111111111111111111111111100011111111111111111111111111110011111111111111111111101111111111111111111101111111111111111111111011111111111111111111111111111111111111111111100000000000000"),
("00000000000000000011111111111111111111111000111111111111111111111111111110011111111011111111111101111111111111111111101111111111111111111111111111111111111101111111111101111111111111111100000000000000"),
("00000000000000000011111111111111111000000011111111111111111101111111111110111111111011111111111101111111111111111111101111111111111111111111111111111111111111111111111111111111111011111100000000000000"),
("00000000000000000011111111111111111000111111111111111111111101111111111110111111111111111111111001111111111111111111001111111111111111111110111111111111111111111111111011111111111011111100000000000000"),
("00000000000000000011111111111111111111111111111111111111111101111111111110111111111111111111111011111111111111111111111111111111111111111110111111111111111111111111111111111111111111111100000000000000"),
("00000000000000000011111111111111110111111111111111111111111111111111111101111111111111111111111011111111111111111111011111111111111111111111111111111111111111111111110111111111110111111000000000000000"),
("00000000000000000111111111111111111111111111111111111111111111111111111101111111111111111111111011111111111111111111011111111111111111111111111111111111111111111111111111111111110111111000000000000000"),
("00000000000000000111111111111111111111111111111111111111111111111111111101111111111111111111111011111111111111111110111111111111111111111111111111111111111111111111101111111111111111111000000000000000"),
("00000000000000000111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111101111111000000000000000"),
("00000000000000000111111111111111101111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111011111111111111111110000000000000000"),
("00000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000011111111111111111111111111111111111111011111111111111110111111111111011111110000000000000000"),
("00000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111011111111111111111111110111111111111111011111111111111101111111111111111111110000000000000000"),
("00000000000000001111111111111111011111111111111111111111111111111111111111111111111110011111111111110111111111111111111111111111000111111111111100101111111111111011111111111110111111100000000000000000"),
("00000000000000001111111111111111011111111111111111111111111111111111111111111111111001011111111111101111111111111111111111111110011011111111111001111111111111110111111111111101111111100000000000000000"),
("00000000000000001111111111111111111111111111111111111111111111111111111110111111110011101111111110011111111101111111110111111100111101111111110011110111111111001111111111111101111111100000000000000000"),
("00000000000000001111111111111111111111111111111111111111111111111111111110011111000111110111111100111111111110111111100111110011111110111111000111111001111100011111111111111011111111000000000000000000"),
("00000000000000001111110000000111111111111111111111111111111111111111111111100000011111110000000011111111111111000000011000000111111111000000011111111100000001111111111111111011111111000000000000000000"),
("00000000000000011111110110011111111111111111111111111111111111111111111111111000111111111100001111111111111111110000111101111111111111110011111111111111110111111111111111110111111110000000000000000000"),
("00000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111110000000000000000000"),
("00000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111100000000000000000000"),
("00000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000"),
("00000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111000000000000000000000"),
("00000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111000000000000000000000"),
("00000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111110000000000000000000000"),
("00000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111100000000000000000000000"),
("00000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111100000000000000000000000"),
("00000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011111111111000000000000000000000000"),
("00000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111110000000000000000000000000"),
("00000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111110000000000000000000000000"),
("00000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111100000000000000000000000000"),
("00000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111111000000000000000000000000000"),
("00000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111110001110001111111111111111111111111111111111111111111111111111110011111111111110000000000000000000000000000"),
("00000000001111111111111111111110000000001111111111111111111111111111111111111111111111100111100101110101110111111111111111111111111111111111111111111111111000111111111111100000000000000000000000000000"),
("00000000001111111111111111110000000010000000000011111111111111111111111111111110111111100111101111110111110111100011111111111111111111111111111111111111110011111111111111000000000000000000000000000000"),
("00000000001111111111111110000111111111111111100000001111111111111111111111100110111111100111101111110111110111101001111111111111111111111111111111111111001111111111111110000000000000000000000000000000"),
("00000000001111111111111000111111111111111111111111100000001111111111111110000110111111111011101111110111110111011111110001111111111111111111111111111100111111111111111110000000000000000000000000000000"),
("00000000011111111111110011111111111111111111111111111111000001111111111110111110111111011011110111110011110111011111110101111111111111111111111111110011111111111111111000000000000000000000000000000000"),
("00000000011111111111001111111111111111111111111111111111111100000111111101111110111111011011110011111001110111011111110111111111111111111111111110001111111111111111110000000000000000000000000000000000"),
("00000000011111111110011111111111111111111111111111111111111111110011111101111110111111011011111101111100110111011111110111111111111111111111110000111111111111111111100000000000000000000000000000000000"),
("00000000011111111100111111111111111111111111111111111111111111111111111101111110111111011011111101111110110111011111110111111111111111111100000111111111111111111111000000000000000000000000000000000000"),
("00000000011111111001111111111111111111111111111111111111111111111111111111111110111110010011111101111110110111011111111011111111111111100000111111111111111111111110000000000000000000000000000000000000"),
("00000000111111111011111111111111111111111111111111111111111111111111111111111110111110000001111101111110110111011111111001111111111000001111111111111111111111111000000000000000000000000000000000000000"),
("00000000111111110111111111111111111111111111111111111111111111111111111111111110111110111101101101110100110111011111111101111111111111111111111111111111111111100000000000000000000000000000000000000000"),
("00000000111111001111111111111111111111111111111111111111111111111111111101111110111110111101100011110001110111101111111110111111111111111111111111111111111111000000000000000000000000000000000000000000"),
("00000000111111111111111111111100000000000000111111111111111111111111111101111110000111111111111111111111111111100101111110111111111111111111111111111111111100000000000000000000000000000000000000000000"),
("00000000011111111111111111110000000000000000000000111111111111111111111101110110011111111111111111111111111111110001111110111111111111111111111111111111110000000000000000000000000000000000000000000000"),
("00000000011111111111111111100000000000000000000000000111111111111111111100001111111111111111111111111111111111111111110100111111111111111111111111111111000000000000000000000000000000000000000000000000"),
("00000000011111111111111110000000000000000000000000000000111111111111111110011111111111111111111111111111111111111111111001111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("00000000011111111111111000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000"),
("00000000001111111111111000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000"),
("00000000001111111111110000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000"),
("00000000000111111111100000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000"),
("00000000000111111111000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000"),
("00000000000011111100000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000110000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000001111111111111111111111111111111000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000001111111111111111111111100000000000000000000000000000011111111111111111111111110000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000011111111111111111111110000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000011111111111111111100000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000011111111111111111000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000011111111111111110000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000001111111111111100000000000000000000000000000000000000000000000001111111111111110000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000000011111111111110000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000001111111111110000000000000000000000000000000000000000000000000000011111111111100000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000111111111110000000000000000000000000000000000000000000000000000001111111111100000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000001111111111000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000011111111000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000111110000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000")
);	

begin

-- Calculate object end boundaries
	objectEndX	<= Draw_Size_X+ObjectStartX;
	objectEndY	<= Draw_Size_Y+ObjectStartY;

-- Signals drawing_X[Y] are active when obects coordinates are being crossed

-- test if ooCoord is in the rectangle defined by Start and End 
	drawing_X	<= '1' when  (oCoord_X  >= ObjectStartX) and  (oCoord_X < objectEndX) else '0';
   drawing_Y	<= '1' when  (oCoord_Y  >= ObjectStartY) and  (oCoord_Y < objectEndY) else '0';

-- calculate offset from start corner 
	bCoord_X 	<= (oCoord_X - ObjectStartX) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 
	bCoord_Y 	<= (oCoord_Y - ObjectStartY) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 
	
	
	process (CLK, resetN)
	begin
		if (resetN = '0') then
			mVGA_RGB	<=  (others => '0') ; 	
			drawing_request	<=  '0' ;
			sig_color <= logo1_Colors;
			sig_mask <= logo1_Mask;

		elsif rising_edge(CLK) then
			
				sig_draw_req <= '0';
				sig_draw_data <= (others => '0');
				
				
				sig_color <= logo1_Colors;
				sig_mask <= logo1_Mask;
					
					
				sig_draw_data <= sig_color(bCoord_Y , bCoord_X);
				sig_draw_req <= sig_mask(bCoord_Y , bCoord_X) and drawing_X and drawing_Y ;
					
			
				mVGA_RGB	<=  sig_draw_data;	 
				drawing_request	<=  sig_draw_req ; 
		
		end if;
	end process;

end architecture;



