library IEEE;
use IEEE.STD_LOGIC_1164.all;
entity logo3 is
port 	(
		
	   CLK  		: in std_logic;
		RESETn		: in std_logic;
		oCoord_X	: in integer;
		oCoord_Y	: in integer;
		ObjectStartX	: in integer;
		ObjectStartY 	: in integer;
		drawing_request	: out std_logic ;
		mVGA_RGB 	: out std_logic_vector(7 downto 0) 
	);
end entity;


architecture behav of logo3 is 

constant object_X_size : integer := 576;
constant object_Y_size : integer := 324;
type ram_array is array(0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic_vector(7 downto 0);
constant object_colors: ram_array := (
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fe",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fd",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fd",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fe",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fe",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fe",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fe",x"fd",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f9",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fa",x"f9",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fe",x"ff",x"ff",x"fe",x"fe",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"f9",x"f9",x"f8",x"f8",x"f8",x"fc",x"fc",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fd",x"fe",x"ff",x"ff",x"ff",x"fe",x"fd",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fa",x"d5",x"d4",x"f4",x"f8",x"f8",x"fc",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fd",x"fe",x"ff",x"ff",x"fe",x"fd",x"fc",x"fc",x"fd",x"fc",x"f8",x"f8",x"f8",x"f9",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"da",x"d5",x"d4",x"d4",x"f4",x"f8",x"f8",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fd",x"fe",x"ff",x"ff",x"fe",x"fd",x"fc",x"fc",x"fd",x"fc",x"f8",x"f8",x"f8",x"f9",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"d6",x"b0",x"b0",x"d4",x"f4",x"f8",x"f8",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fd",x"fe",x"ff",x"ff",x"fe",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f9",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"b5",x"90",x"b0",x"b4",x"d4",x"f4",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fd",x"fe",x"ff",x"ff",x"fe",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f9",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"b5",x"8c",x"90",x"b0",x"d4",x"d4",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fd",x"fe",x"ff",x"ff",x"fe",x"fd",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"fa",x"f6",x"f6",x"f6",x"d2",x"d2",x"d2",x"d2",x"ce",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"cd",x"ce",x"ce",x"d2",x"f2",x"f2",x"f6",x"f6",x"fb",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"da",x"b1",x"8c",x"90",x"b0",x"d4",x"d4",x"d4",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fd",x"fe",x"ff",x"ff",x"fe",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"da",x"d6",x"d2",x"d2",x"cd",x"cd",x"cd",x"a9",x"a9",x"a9",x"a9",x"85",x"85",x"84",x"84",x"60",x"60",x"60",x"80",x"80",x"84",x"84",x"84",x"84",x"a5",x"a5",x"a9",x"a9",x"a9",x"cd",x"ce",x"d2",x"d2",x"d6",x"d6",x"db",x"fb",x"ff",x"da",x"d5",x"90",x"8c",x"90",x"b0",x"b4",x"d4",x"d4",x"f4",x"f8",x"fd",x"fd",x"fe",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fe",x"fe",x"ff",x"fe",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f9",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"da",x"d6",x"d6",x"d2",x"ad",x"a9",x"a5",x"a4",x"a4",x"84",x"80",x"80",x"60",x"60",x"60",x"64",x"64",x"64",x"64",x"64",x"64",x"64",x"64",x"64",x"64",x"64",x"64",x"64",x"64",x"64",x"44",x"44",x"44",x"44",x"40",x"40",x"40",x"60",x"64",x"64",x"85",x"85",x"a9",x"a9",x"c9",x"ad",x"8d",x"8c",x"8c",x"8c",x"90",x"b4",x"d4",x"d4",x"f8",x"f8",x"fd",x"fd",x"fe",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fd",x"fe",x"ff",x"ff",x"fe",x"fd",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f9",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fa",x"d6",x"d6",x"b2",x"ad",x"a9",x"89",x"84",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"64",x"64",x"64",x"68",x"69",x"69",x"69",x"69",x"89",x"8d",x"8d",x"8d",x"89",x"89",x"89",x"69",x"69",x"69",x"68",x"48",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"84",x"88",x"8c",x"8c",x"8c",x"90",x"b0",x"d4",x"d4",x"f4",x"f8",x"f9",x"fd",x"fe",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fd",x"fe",x"ff",x"ff",x"fe",x"fd",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"d2",x"cd",x"a9",x"a4",x"84",x"60",x"60",x"60",x"64",x"84",x"89",x"89",x"8d",x"ad",x"b1",x"d2",x"d2",x"d6",x"d6",x"d6",x"d6",x"d6",x"d6",x"d6",x"d6",x"d6",x"d6",x"d6",x"d2",x"d2",x"d2",x"d2",x"d2",x"d2",x"d2",x"ce",x"cd",x"cd",x"cd",x"a9",x"a9",x"a9",x"89",x"89",x"68",x"64",x"44",x"20",x"20",x"00",x"44",x"68",x"8c",x"8c",x"8c",x"8c",x"b0",x"d4",x"d4",x"f4",x"f8",x"f9",x"fd",x"fe",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fd",x"fe",x"ff",x"ff",x"fe",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"d9",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"d6",x"d2",x"ad",x"a9",x"84",x"80",x"80",x"60",x"60",x"85",x"85",x"89",x"8d",x"92",x"b2",x"b6",x"b6",x"da",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fb",x"fa",x"f6",x"f6",x"f6",x"f6",x"f6",x"f6",x"f2",x"f2",x"f2",x"f2",x"f2",x"f2",x"ee",x"ee",x"ee",x"ed",x"ed",x"cd",x"cd",x"ad",x"ad",x"89",x"68",x"44",x"24",x"20",x"44",x"84",x"8c",x"ac",x"8c",x"8c",x"b0",x"b0",x"d4",x"d4",x"f8",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fd",x"fe",x"ff",x"fe",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"d9",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"d2",x"a9",x"a5",x"84",x"60",x"60",x"60",x"64",x"68",x"89",x"b2",x"d6",x"d6",x"d6",x"db",x"db",x"df",x"df",x"df",x"db",x"db",x"fa",x"fa",x"f6",x"f6",x"f6",x"f2",x"f2",x"f2",x"f2",x"f2",x"ee",x"ed",x"ed",x"ed",x"ed",x"ed",x"ed",x"ed",x"ed",x"ed",x"ed",x"ed",x"ed",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"c9",x"c9",x"c9",x"c9",x"a8",x"88",x"ac",x"ac",x"ac",x"8c",x"b0",x"b0",x"d0",x"d4",x"f4",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fd",x"fe",x"fe",x"fe",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"f6",x"d6",x"d2",x"ad",x"a5",x"80",x"60",x"60",x"60",x"64",x"89",x"8d",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"fa",x"f6",x"f6",x"f2",x"f2",x"f2",x"ed",x"ed",x"ed",x"ed",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e5",x"e5",x"e5",x"e5",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"a8",x"ac",x"ac",x"ac",x"8c",x"b0",x"b0",x"d0",x"d4",x"f4",x"f8",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fe",x"fe",x"fe",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"d9",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"db",x"d2",x"a9",x"a4",x"80",x"60",x"60",x"60",x"60",x"68",x"8d",x"b2",x"d6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"f6",x"f6",x"f2",x"f2",x"ee",x"ed",x"ed",x"ed",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e5",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e5",x"e9",x"e9",x"a8",x"a8",x"ac",x"ac",x"b0",x"b0",x"b0",x"d0",x"d4",x"f4",x"f8",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fd",x"fc",x"fc",x"fd",x"fe",x"fe",x"fe",x"fe",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"d9",x"da",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"d6",x"d2",x"b2",x"ad",x"89",x"80",x"60",x"60",x"60",x"64",x"69",x"8d",x"b1",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"f6",x"f2",x"f2",x"ed",x"ed",x"e9",x"e9",x"e9",x"e5",x"e5",x"e4",x"e4",x"c4",x"c4",x"e4",x"e4",x"c4",x"c4",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c4",x"c4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"c8",x"a8",x"a8",x"ac",x"b0",x"b0",x"b0",x"b0",x"d4",x"f4",x"f8",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fd",x"fd",x"fe",x"fe",x"fe",x"fd",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"d8",x"d9",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"d2",x"a9",x"84",x"60",x"60",x"60",x"60",x"40",x"65",x"89",x"b2",x"d6",x"db",x"ff",x"ff",x"ff",x"fb",x"fb",x"fa",x"f6",x"f6",x"f6",x"f2",x"ed",x"ed",x"e9",x"e9",x"e9",x"e5",x"e5",x"e4",x"e4",x"e4",x"c4",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"e0",x"e4",x"e4",x"c4",x"a4",x"a8",x"ac",x"b0",x"90",x"b0",x"b0",x"d0",x"f4",x"f4",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fd",x"fd",x"fe",x"fe",x"fe",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"fc",x"f8",x"d8",x"d9",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"d2",x"ce",x"a9",x"a5",x"80",x"60",x"60",x"64",x"64",x"89",x"8d",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"f6",x"f2",x"f2",x"ed",x"ed",x"e9",x"e4",x"e4",x"e4",x"e4",x"c4",x"c4",x"c4",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"c0",x"a0",x"a0",x"a4",x"a8",x"ac",x"90",x"90",x"90",x"b0",x"d0",x"f4",x"f4",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fd",x"fd",x"fe",x"fe",x"fe",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"d8",x"d8",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"d2",x"ad",x"a9",x"84",x"60",x"60",x"60",x"60",x"85",x"8d",x"b2",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"f6",x"f6",x"f2",x"f2",x"ee",x"ed",x"e9",x"e5",x"e5",x"e4",x"c4",x"c4",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"88",x"8c",x"90",x"90",x"90",x"b0",x"d0",x"d4",x"f4",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fd",x"fe",x"fe",x"fe",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"d8",x"d8",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"d6",x"d2",x"cd",x"ad",x"a9",x"84",x"84",x"64",x"64",x"64",x"89",x"8d",x"b2",x"d6",x"db",x"fb",x"fb",x"ff",x"ff",x"fb",x"fa",x"f6",x"f2",x"f2",x"ed",x"ed",x"e9",x"e9",x"e5",x"c4",x"c4",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"80",x"80",x"88",x"8c",x"90",x"90",x"90",x"b0",x"d0",x"d4",x"f4",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fe",x"fe",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f9",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d2",x"cd",x"c9",x"a4",x"60",x"60",x"60",x"64",x"68",x"8d",x"91",x"b6",x"da",x"fb",x"ff",x"fb",x"fb",x"fb",x"f7",x"f6",x"f6",x"f2",x"f2",x"ed",x"e9",x"e9",x"e5",x"e5",x"e4",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"88",x"ac",x"90",x"90",x"90",x"b0",x"b0",x"d4",x"f4",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fd",x"fd",x"fe",x"fe",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"d5",x"da",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"d6",x"d6",x"b2",x"ad",x"a9",x"85",x"84",x"84",x"64",x"84",x"89",x"8d",x"b2",x"b6",x"d6",x"fb",x"fb",x"ff",x"fb",x"fb",x"f6",x"f6",x"f2",x"f2",x"ed",x"ed",x"e9",x"e9",x"e5",x"e4",x"c4",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"64",x"64",x"64",x"64",x"64",x"84",x"84",x"85",x"85",x"85",x"89",x"89",x"85",x"85",x"85",x"85",x"85",x"89",x"89",x"89",x"89",x"69",x"65",x"65",x"65",x"65",x"65",x"64",x"64",x"64",x"64",x"64",x"60",x"60",x"60",x"60",x"80",x"80",x"84",x"88",x"8c",x"8c",x"90",x"b0",x"b0",x"d4",x"f4",x"f4",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fd",x"fd",x"fe",x"fe",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"d4",x"d9",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"d6",x"ce",x"a9",x"85",x"80",x"60",x"60",x"64",x"64",x"69",x"b2",x"b6",x"d6",x"db",x"fb",x"fb",x"fb",x"fb",x"fa",x"f6",x"f6",x"f2",x"f1",x"ed",x"ed",x"e9",x"e9",x"e5",x"e4",x"c4",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"64",x"64",x"44",x"64",x"68",x"68",x"68",x"89",x"89",x"a9",x"a9",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"8d",x"8d",x"8d",x"89",x"89",x"69",x"69",x"69",x"69",x"65",x"64",x"44",x"44",x"60",x"80",x"80",x"64",x"68",x"6c",x"8c",x"90",x"b0",x"b0",x"d4",x"d4",x"f4",x"f8",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fd",x"fe",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"d8",x"d9",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"d6",x"d2",x"ae",x"a9",x"a9",x"85",x"84",x"84",x"84",x"85",x"89",x"8d",x"91",x"b6",x"db",x"fb",x"fb",x"fb",x"fb",x"fa",x"f6",x"f6",x"f2",x"f2",x"f1",x"ed",x"e9",x"e9",x"e8",x"c4",x"c4",x"c4",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"64",x"84",x"88",x"88",x"88",x"89",x"89",x"89",x"a9",x"a9",x"a9",x"a9",x"c9",x"c9",x"c9",x"c9",x"c9",x"c9",x"c9",x"c9",x"c9",x"c9",x"c9",x"c9",x"c9",x"e9",x"cd",x"cd",x"cd",x"cd",x"cd",x"c9",x"c9",x"c9",x"a9",x"a9",x"a9",x"a9",x"a9",x"89",x"89",x"89",x"84",x"84",x"64",x"64",x"68",x"6c",x"6c",x"90",x"90",x"b0",x"d4",x"d4",x"f4",x"f8",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"d8",x"d9",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fa",x"d6",x"ae",x"a9",x"85",x"80",x"60",x"60",x"60",x"64",x"89",x"8d",x"b2",x"d6",x"da",x"fb",x"fb",x"fb",x"fb",x"fb",x"f6",x"f6",x"f2",x"ed",x"ed",x"ed",x"ed",x"e9",x"e9",x"e4",x"e4",x"c0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"60",x"44",x"64",x"64",x"88",x"89",x"ad",x"ad",x"cd",x"cd",x"cd",x"c9",x"e9",x"e9",x"e9",x"e9",x"e8",x"e8",x"e8",x"e8",x"e4",x"c4",x"c4",x"c4",x"c4",x"c4",x"c4",x"c4",x"e4",x"e9",x"e5",x"e4",x"e4",x"e4",x"e4",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"c9",x"c9",x"c9",x"c9",x"a9",x"88",x"68",x"68",x"6c",x"6c",x"70",x"90",x"90",x"b0",x"b4",x"d4",x"d4",x"f8",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"d8",x"d8",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"d2",x"ad",x"a9",x"89",x"85",x"85",x"64",x"64",x"65",x"89",x"89",x"ad",x"d2",x"d6",x"d6",x"fa",x"fb",x"fb",x"f6",x"f6",x"f6",x"f2",x"f2",x"ed",x"e9",x"e9",x"e5",x"e5",x"e4",x"c4",x"c4",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"60",x"60",x"60",x"60",x"60",x"64",x"64",x"64",x"84",x"84",x"a8",x"a9",x"a9",x"c9",x"c9",x"c9",x"e9",x"e9",x"c9",x"c5",x"c5",x"c4",x"c4",x"a4",x"84",x"84",x"84",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"84",x"a4",x"a4",x"a4",x"c4",x"c4",x"c4",x"c4",x"e4",x"e9",x"e9",x"e9",x"c9",x"a9",x"a9",x"8d",x"8c",x"8c",x"90",x"90",x"90",x"b0",x"d4",x"d4",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"d4",x"d5",x"d6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"d2",x"ad",x"85",x"60",x"60",x"60",x"60",x"64",x"89",x"8d",x"92",x"b6",x"d6",x"fb",x"fb",x"fb",x"fb",x"f6",x"f6",x"f2",x"f1",x"ed",x"e9",x"e9",x"e9",x"e9",x"e5",x"e4",x"e0",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"60",x"60",x"64",x"64",x"64",x"64",x"68",x"68",x"a9",x"c9",x"c9",x"c9",x"e9",x"e9",x"e5",x"e5",x"e5",x"c4",x"c0",x"a0",x"a0",x"a0",x"80",x"60",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"40",x"40",x"60",x"60",x"80",x"a0",x"a0",x"c0",x"c4",x"e4",x"e5",x"e9",x"c9",x"c9",x"c9",x"ad",x"ac",x"ac",x"8c",x"8c",x"b0",x"d4",x"d4",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"d4",x"b0",x"b1",x"d6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"d2",x"ae",x"ad",x"89",x"84",x"64",x"64",x"64",x"64",x"89",x"8d",x"ad",x"b2",x"d6",x"d6",x"f6",x"f6",x"f6",x"f6",x"f6",x"f2",x"f2",x"ed",x"ed",x"e9",x"e4",x"e4",x"e4",x"e4",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"64",x"64",x"88",x"89",x"89",x"a9",x"a9",x"a9",x"a9",x"c9",x"c5",x"c5",x"c4",x"a4",x"a4",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"40",x"44",x"44",x"44",x"48",x"68",x"68",x"68",x"64",x"64",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"a0",x"c0",x"c4",x"c4",x"c5",x"c8",x"ac",x"ac",x"ac",x"ac",x"b0",x"d4",x"d4",x"d8",x"f8",x"fc",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fe",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"fc",x"fc",x"f8",x"f8",x"b0",x"8c",x"89",x"8d",x"d6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"d2",x"ad",x"85",x"84",x"60",x"60",x"60",x"60",x"64",x"89",x"ad",x"b2",x"d6",x"f6",x"fa",x"f6",x"f6",x"f6",x"f2",x"f2",x"ed",x"ed",x"e9",x"e9",x"e9",x"e5",x"e4",x"e4",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"64",x"64",x"64",x"88",x"89",x"ad",x"cd",x"cd",x"e9",x"e9",x"e9",x"c5",x"a4",x"a4",x"80",x"80",x"60",x"60",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"64",x"88",x"a8",x"ac",x"d0",x"d0",x"d0",x"d4",x"d0",x"d0",x"ac",x"a8",x"88",x"64",x"40",x"40",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"40",x"80",x"80",x"80",x"80",x"a8",x"a8",x"ac",x"ac",x"b0",x"b0",x"b4",x"d4",x"d4",x"d8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fe",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"fc",x"fd",x"f8",x"d4",x"8c",x"44",x"44",x"8d",x"d6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"db",x"d7",x"d2",x"cd",x"a9",x"85",x"64",x"60",x"60",x"64",x"64",x"89",x"89",x"ad",x"b2",x"d6",x"d6",x"f6",x"f6",x"f6",x"f2",x"f2",x"f2",x"f2",x"ed",x"ed",x"e9",x"e9",x"e4",x"e4",x"c4",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"64",x"64",x"64",x"89",x"89",x"a9",x"c9",x"c9",x"c9",x"e9",x"e9",x"c9",x"c4",x"c4",x"a4",x"80",x"80",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"60",x"60",x"84",x"88",x"ac",x"d0",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"d4",x"d0",x"ac",x"88",x"64",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"20",x"40",x"64",x"68",x"8c",x"90",x"90",x"b0",x"b0",x"d4",x"d4",x"f4",x"f8",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fe",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"b0",x"44",x"40",x"64",x"89",x"d2",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"d6",x"b2",x"ae",x"a5",x"a0",x"80",x"60",x"40",x"40",x"64",x"89",x"ad",x"b2",x"d2",x"d6",x"f6",x"fb",x"fb",x"f6",x"f2",x"ee",x"ed",x"ed",x"e9",x"e9",x"e9",x"e9",x"e5",x"e4",x"c4",x"c0",x"c0",x"a0",x"80",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"64",x"64",x"48",x"68",x"89",x"a9",x"cd",x"e9",x"e9",x"e9",x"e5",x"e5",x"c4",x"c0",x"a0",x"80",x"60",x"60",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"64",x"88",x"ac",x"d0",x"f9",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"f8",x"d4",x"ac",x"88",x"64",x"40",x"40",x"40",x"40",x"20",x"00",x"00",x"00",x"00",x"24",x"48",x"6c",x"70",x"90",x"b0",x"b0",x"d4",x"f4",x"f4",x"f8",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fe",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"d0",x"68",x"40",x"40",x"44",x"89",x"b2",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"d2",x"ad",x"a9",x"85",x"84",x"64",x"60",x"64",x"64",x"89",x"89",x"ad",x"b1",x"d2",x"d2",x"f2",x"f2",x"f2",x"f2",x"f2",x"f2",x"ed",x"ed",x"e9",x"e9",x"e9",x"e4",x"e4",x"e4",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"60",x"60",x"64",x"64",x"64",x"64",x"64",x"88",x"88",x"a9",x"a9",x"c9",x"c9",x"c9",x"c9",x"c5",x"c4",x"c4",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"68",x"ac",x"d4",x"d8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"d4",x"ac",x"64",x"40",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"40",x"68",x"8c",x"90",x"90",x"90",x"b0",x"d4",x"f4",x"f4",x"f8",x"fc",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"fc",x"f8",x"f8",x"f4",x"8c",x"44",x"00",x"00",x"40",x"85",x"cd",x"f6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"d2",x"ad",x"89",x"84",x"60",x"60",x"60",x"60",x"64",x"69",x"8d",x"ad",x"d2",x"f6",x"f6",x"f6",x"f6",x"f2",x"f2",x"ed",x"ed",x"e9",x"e9",x"e9",x"e9",x"e5",x"e4",x"e4",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"64",x"64",x"64",x"64",x"68",x"68",x"89",x"a9",x"a9",x"c9",x"e9",x"e9",x"e9",x"e5",x"c4",x"a0",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"44",x"68",x"b0",x"d4",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"d4",x"ac",x"64",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"84",x"8c",x"90",x"90",x"90",x"b0",x"d4",x"d4",x"f4",x"f8",x"f8",x"fc",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f4",x"b0",x"68",x"00",x"00",x"20",x"40",x"80",x"cd",x"f7",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"d6",x"d2",x"cd",x"a9",x"85",x"84",x"64",x"64",x"64",x"64",x"68",x"89",x"8d",x"ad",x"d2",x"d2",x"d2",x"f2",x"f2",x"f2",x"f2",x"ee",x"ed",x"ed",x"e9",x"e9",x"e5",x"e4",x"e4",x"e4",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"64",x"64",x"64",x"68",x"89",x"ad",x"cd",x"cd",x"c9",x"e9",x"e9",x"c5",x"c4",x"a4",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"64",x"8c",x"d0",x"d4",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"d4",x"ac",x"64",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"84",x"8c",x"8c",x"90",x"90",x"b0",x"b4",x"d4",x"f4",x"f4",x"f8",x"fc",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"fc",x"fc",x"fc",x"f8",x"d4",x"8c",x"40",x"20",x"20",x"20",x"40",x"64",x"a9",x"d6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"b2",x"ad",x"89",x"80",x"60",x"60",x"60",x"60",x"64",x"68",x"8d",x"ad",x"b1",x"d2",x"f6",x"f2",x"f2",x"f2",x"ed",x"ed",x"ed",x"e9",x"e9",x"e9",x"e9",x"e5",x"e4",x"c4",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"64",x"64",x"64",x"64",x"64",x"68",x"88",x"a9",x"c9",x"ed",x"ed",x"e9",x"e9",x"e5",x"c5",x"a0",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"20",x"20",x"40",x"64",x"8c",x"d4",x"f9",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fd",x"f9",x"d5",x"ac",x"64",x"40",x"40",x"40",x"40",x"40",x"40",x"64",x"8c",x"8c",x"90",x"90",x"b0",x"b0",x"d0",x"d4",x"f4",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"fc",x"f8",x"f4",x"cc",x"80",x"60",x"40",x"20",x"00",x"20",x"60",x"ad",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"f2",x"c9",x"a9",x"85",x"64",x"64",x"44",x"44",x"64",x"64",x"89",x"a9",x"cd",x"cd",x"d2",x"d2",x"d2",x"f2",x"f2",x"f1",x"ed",x"ed",x"e9",x"e9",x"e5",x"e5",x"e5",x"e4",x"e4",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"40",x"44",x"44",x"64",x"88",x"89",x"a9",x"a9",x"cd",x"e9",x"e9",x"e9",x"e5",x"c4",x"c0",x"a0",x"80",x"64",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"68",x"b0",x"d4",x"f8",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"f9",x"d4",x"ac",x"64",x"40",x"40",x"40",x"40",x"40",x"64",x"88",x"8c",x"8c",x"90",x"b0",x"b0",x"b0",x"d4",x"d4",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"fc",x"f8",x"f8",x"ec",x"c4",x"a0",x"60",x"20",x"00",x"00",x"40",x"64",x"a8",x"f2",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"f6",x"d6",x"d2",x"cd",x"a5",x"80",x"80",x"60",x"60",x"60",x"64",x"64",x"69",x"8d",x"cd",x"ee",x"f2",x"f2",x"f2",x"f2",x"f1",x"ed",x"ed",x"e9",x"e9",x"e5",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"64",x"64",x"64",x"64",x"64",x"64",x"68",x"a9",x"a9",x"c9",x"ed",x"e9",x"e9",x"e5",x"e5",x"c0",x"a0",x"80",x"60",x"40",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"20",x"20",x"00",x"20",x"48",x"8c",x"d8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fe",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fe",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"f8",x"d4",x"8c",x"40",x"40",x"40",x"40",x"40",x"64",x"88",x"8c",x"8c",x"b0",x"b0",x"b0",x"b0",x"d4",x"d4",x"f8",x"f8",x"f9",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f0",x"e4",x"c0",x"a0",x"40",x"20",x"00",x"20",x"40",x"60",x"a9",x"f2",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"f7",x"d2",x"a9",x"a5",x"84",x"84",x"64",x"40",x"20",x"40",x"64",x"89",x"a9",x"ad",x"cd",x"cd",x"ee",x"ed",x"ed",x"ed",x"ed",x"e9",x"e9",x"e9",x"e5",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"44",x"44",x"44",x"68",x"89",x"a9",x"cd",x"cd",x"ed",x"e9",x"e9",x"e9",x"c5",x"a4",x"a0",x"80",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"40",x"20",x"20",x"00",x"00",x"20",x"44",x"90",x"d4",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fe",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"fc",x"f8",x"b0",x"68",x"40",x"40",x"20",x"40",x"64",x"88",x"8c",x"ac",x"b0",x"b0",x"b0",x"b0",x"d4",x"d4",x"f8",x"f8",x"f9",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f0",x"e8",x"e4",x"c0",x"a0",x"80",x"20",x"00",x"20",x"40",x"60",x"84",x"d2",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"f6",x"d2",x"cd",x"a5",x"80",x"60",x"60",x"60",x"64",x"44",x"44",x"48",x"89",x"ad",x"cd",x"ed",x"ee",x"ee",x"ed",x"ed",x"ed",x"e9",x"e9",x"e5",x"e4",x"e4",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"64",x"64",x"64",x"68",x"69",x"89",x"a9",x"c9",x"ed",x"ed",x"e9",x"e9",x"c5",x"c4",x"a0",x"80",x"60",x"40",x"40",x"20",x"20",x"40",x"40",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"00",x"00",x"00",x"20",x"20",x"20",x"00",x"00",x"00",x"44",x"6c",x"d4",x"f9",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fe",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fe",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"fc",x"fc",x"d4",x"8c",x"64",x"20",x"20",x"20",x"40",x"64",x"8c",x"b0",x"b0",x"b0",x"b0",x"b0",x"b4",x"d4",x"f8",x"f8",x"f9",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"d4",x"cc",x"c8",x"e0",x"c0",x"c0",x"60",x"00",x"00",x"20",x"40",x"60",x"89",x"d6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f7",x"d2",x"a9",x"85",x"84",x"64",x"60",x"40",x"40",x"40",x"64",x"88",x"ad",x"ad",x"cd",x"cd",x"ed",x"ed",x"ed",x"ed",x"e9",x"e9",x"e9",x"e5",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"64",x"44",x"44",x"44",x"68",x"89",x"a9",x"c9",x"c9",x"e9",x"e9",x"e9",x"e5",x"c4",x"a0",x"80",x"80",x"60",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"20",x"20",x"20",x"00",x"00",x"00",x"20",x"68",x"b0",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fe",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"fc",x"f8",x"b0",x"68",x"20",x"20",x"20",x"40",x"44",x"8c",x"b0",x"b0",x"b0",x"b0",x"b0",x"b4",x"d4",x"f8",x"f8",x"f9",x"f9",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"d4",x"d0",x"c8",x"c0",x"e0",x"e0",x"a0",x"80",x"20",x"00",x"00",x"20",x"60",x"84",x"f6",x"ff",x"ff",x"ff",x"df",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"f6",x"d2",x"ad",x"89",x"60",x"60",x"40",x"40",x"40",x"60",x"64",x"64",x"89",x"ad",x"cd",x"ed",x"ee",x"ed",x"ed",x"e9",x"e9",x"e9",x"e9",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"64",x"64",x"68",x"48",x"68",x"69",x"89",x"a9",x"c9",x"e9",x"e9",x"e9",x"e5",x"c5",x"c0",x"a0",x"80",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"44",x"8c",x"d4",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fe",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fe",x"fd",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f8",x"d4",x"88",x"40",x"20",x"20",x"20",x"44",x"68",x"b0",x"b0",x"b0",x"b0",x"b0",x"b4",x"d4",x"d4",x"f8",x"f9",x"f9",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"d4",x"ac",x"a0",x"c0",x"c0",x"e0",x"c0",x"60",x"00",x"00",x"00",x"20",x"60",x"a9",x"f6",x"ff",x"ff",x"df",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"d2",x"ad",x"a9",x"84",x"80",x"60",x"40",x"40",x"40",x"40",x"64",x"a9",x"c9",x"cd",x"ed",x"ed",x"ed",x"ed",x"e9",x"e9",x"e9",x"e4",x"e4",x"e5",x"e5",x"e5",x"e4",x"e4",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"44",x"44",x"68",x"69",x"8d",x"ad",x"cd",x"e9",x"e9",x"e9",x"e5",x"c4",x"a0",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"64",x"88",x"b0",x"d4",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fe",x"fe",x"ff",x"ff",x"ff",x"fe",x"fe",x"fe",x"fd",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f4",x"8c",x"44",x"20",x"00",x"00",x"20",x"68",x"8c",x"8c",x"b0",x"b0",x"b0",x"b4",x"d4",x"d4",x"f8",x"f9",x"f9",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"d4",x"ac",x"a4",x"a0",x"a0",x"c0",x"e0",x"a0",x"60",x"00",x"00",x"20",x"40",x"60",x"a8",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"f6",x"d6",x"d2",x"ad",x"89",x"84",x"60",x"60",x"40",x"60",x"60",x"60",x"64",x"84",x"a9",x"cd",x"ed",x"ed",x"ed",x"e9",x"e9",x"e9",x"e9",x"e5",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"64",x"64",x"64",x"64",x"64",x"64",x"84",x"89",x"89",x"a9",x"c9",x"e9",x"e9",x"e9",x"e5",x"c5",x"c0",x"a0",x"80",x"60",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"68",x"ac",x"b0",x"d4",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fe",x"fe",x"ff",x"ff",x"ff",x"fe",x"fe",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fc",x"fc",x"f8",x"f8",x"f8",x"b0",x"64",x"20",x"00",x"00",x"00",x"48",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"d4",x"d4",x"f8",x"f9",x"f9",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"f8",x"f8",x"f4",x"d0",x"88",x"84",x"80",x"c0",x"e0",x"c0",x"a0",x"40",x"20",x"20",x"20",x"40",x"60",x"ad",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"f6",x"d2",x"cd",x"a5",x"84",x"60",x"60",x"60",x"40",x"40",x"44",x"44",x"88",x"c9",x"c9",x"c9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e5",x"e5",x"e5",x"e4",x"e0",x"e0",x"e4",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"44",x"44",x"64",x"89",x"a9",x"cd",x"c9",x"e9",x"e9",x"e9",x"e5",x"c4",x"a4",x"a0",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"88",x"b0",x"d4",x"d4",x"f8",x"f8",x"f8",x"f9",x"fd",x"fe",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fd",x"fd",x"fd",x"fe",x"fe",x"ff",x"ff",x"ff",x"ff",x"fe",x"fe",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"b0",x"68",x"24",x"00",x"00",x"00",x"44",x"6c",x"8c",x"90",x"b0",x"b0",x"b0",x"d4",x"d4",x"f4",x"f9",x"f9",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"fc",x"f8",x"f8",x"f8",x"f9",x"d4",x"ac",x"84",x"80",x"80",x"a0",x"c0",x"e0",x"a0",x"60",x"20",x"00",x"20",x"40",x"60",x"a9",x"f7",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"f6",x"d6",x"d2",x"ad",x"a9",x"84",x"60",x"60",x"60",x"60",x"60",x"84",x"84",x"84",x"88",x"c9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e5",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"80",x"60",x"64",x"64",x"64",x"64",x"64",x"84",x"88",x"a9",x"a9",x"c9",x"e9",x"e9",x"e9",x"e5",x"c4",x"c0",x"a0",x"80",x"80",x"60",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"64",x"88",x"b0",x"d4",x"d4",x"f8",x"f8",x"f8",x"fd",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fd",x"fd",x"fe",x"fe",x"ff",x"ff",x"ff",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"d4",x"8c",x"24",x"00",x"00",x"00",x"24",x"68",x"8c",x"b0",x"b0",x"b0",x"b0",x"d4",x"d4",x"f4",x"f9",x"f9",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"fc",x"f8",x"f8",x"f8",x"f9",x"f4",x"b0",x"88",x"80",x"80",x"80",x"a0",x"e0",x"c0",x"a0",x"60",x"20",x"00",x"20",x"20",x"64",x"ce",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"db",x"d6",x"ae",x"a5",x"80",x"80",x"60",x"40",x"40",x"40",x"44",x"64",x"88",x"a9",x"c9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e5",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"44",x"44",x"68",x"89",x"a9",x"c9",x"c9",x"e9",x"e9",x"e9",x"e5",x"c4",x"a4",x"a0",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"40",x"40",x"40",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"60",x"60",x"60",x"60",x"84",x"88",x"ac",x"b0",x"d0",x"d4",x"f8",x"f8",x"f8",x"fd",x"fe",x"fe",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fe",x"fe",x"ff",x"ff",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"d4",x"8c",x"44",x"00",x"00",x"00",x"24",x"48",x"8c",x"b0",x"b0",x"b0",x"b0",x"d0",x"d4",x"f4",x"f9",x"f9",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"fc",x"f8",x"f8",x"f8",x"f9",x"f5",x"b0",x"88",x"80",x"80",x"80",x"80",x"a0",x"c0",x"c0",x"a0",x"60",x"20",x"00",x"00",x"40",x"84",x"cd",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"f7",x"d6",x"d2",x"ad",x"89",x"65",x"60",x"60",x"60",x"60",x"60",x"60",x"84",x"84",x"a8",x"c9",x"c9",x"e9",x"e9",x"e9",x"e5",x"e5",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"64",x"64",x"64",x"64",x"85",x"89",x"a9",x"a9",x"c9",x"c9",x"e9",x"e9",x"c5",x"c4",x"c4",x"a0",x"80",x"60",x"60",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"a8",x"ac",x"b0",x"b0",x"d4",x"f4",x"f8",x"f8",x"fd",x"fd",x"fe",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f4",x"b0",x"48",x"00",x"00",x"00",x"24",x"48",x"8c",x"b0",x"b0",x"b0",x"b0",x"d0",x"d4",x"d4",x"f8",x"f9",x"f9",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"ac",x"80",x"80",x"80",x"80",x"80",x"a0",x"c0",x"c0",x"a0",x"40",x"00",x"00",x"20",x"60",x"a5",x"f6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f2",x"ce",x"a9",x"a5",x"80",x"60",x"40",x"40",x"60",x"60",x"84",x"84",x"a4",x"c5",x"e9",x"e9",x"e9",x"e5",x"e5",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"44",x"44",x"44",x"64",x"88",x"a9",x"c9",x"c9",x"e9",x"e9",x"e5",x"c5",x"c4",x"a4",x"a0",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"84",x"88",x"8c",x"b0",x"b0",x"d4",x"f4",x"f8",x"f8",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f4",x"d0",x"68",x"20",x"00",x"00",x"20",x"44",x"6c",x"90",x"90",x"b0",x"b0",x"b0",x"d4",x"d4",x"f4",x"f8",x"f9",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f4",x"b0",x"84",x"80",x"80",x"60",x"60",x"80",x"a0",x"e0",x"e0",x"80",x"40",x"00",x"00",x"20",x"60",x"c9",x"f6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f7",x"d2",x"d2",x"ad",x"89",x"84",x"60",x"60",x"60",x"60",x"60",x"60",x"84",x"a4",x"a4",x"c4",x"c4",x"e5",x"e5",x"e5",x"e5",x"e5",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"44",x"64",x"64",x"88",x"88",x"a9",x"c9",x"c9",x"c9",x"e9",x"e4",x"c4",x"c4",x"a0",x"a0",x"80",x"80",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"00",x"20",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a4",x"88",x"8c",x"b0",x"b0",x"b0",x"d4",x"f4",x"f8",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"68",x"20",x"20",x"20",x"20",x"24",x"6c",x"90",x"90",x"90",x"b0",x"b0",x"d4",x"d4",x"d4",x"f8",x"f8",x"f9",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"d0",x"88",x"80",x"80",x"60",x"60",x"60",x"80",x"c0",x"e0",x"a0",x"60",x"20",x"00",x"20",x"40",x"84",x"cd",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"ce",x"a9",x"84",x"60",x"40",x"40",x"20",x"40",x"40",x"64",x"84",x"a4",x"c9",x"c9",x"e9",x"e9",x"e5",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"64",x"44",x"44",x"44",x"44",x"64",x"88",x"a9",x"c9",x"e9",x"e9",x"e5",x"e5",x"c5",x"c4",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"60",x"80",x"80",x"60",x"60",x"80",x"80",x"a0",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a4",x"a8",x"ac",x"b0",x"b0",x"b0",x"d4",x"f4",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"88",x"40",x"20",x"20",x"00",x"20",x"68",x"90",x"8c",x"8c",x"b0",x"b0",x"d0",x"d4",x"d4",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"d0",x"a8",x"84",x"60",x"80",x"80",x"60",x"60",x"a0",x"c0",x"c0",x"a0",x"40",x"20",x"20",x"20",x"40",x"65",x"d2",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"d6",x"d6",x"d2",x"cd",x"a9",x"84",x"60",x"60",x"40",x"40",x"60",x"60",x"80",x"80",x"a4",x"c4",x"c4",x"e5",x"e5",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"64",x"64",x"64",x"64",x"84",x"88",x"a9",x"a9",x"c9",x"c9",x"e5",x"c5",x"c4",x"a4",x"a4",x"a0",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"a4",x"a8",x"ac",x"b0",x"b0",x"b0",x"d4",x"d4",x"f4",x"f8",x"f9",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"8c",x"44",x"20",x"20",x"00",x"20",x"68",x"8c",x"8c",x"8c",x"b0",x"b0",x"d0",x"d4",x"d4",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"d0",x"cc",x"84",x"60",x"80",x"80",x"60",x"60",x"80",x"a0",x"a0",x"a0",x"80",x"60",x"20",x"00",x"00",x"40",x"a9",x"f2",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"ce",x"a9",x"a5",x"80",x"80",x"60",x"60",x"40",x"40",x"64",x"84",x"a4",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"44",x"44",x"48",x"68",x"88",x"a9",x"c9",x"e9",x"e9",x"e9",x"e5",x"e5",x"c0",x"a0",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"20",x"20",x"40",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"80",x"a0",x"c0",x"c0",x"a0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"a4",x"a8",x"ac",x"b0",x"b0",x"b0",x"b0",x"d4",x"d4",x"f8",x"f9",x"f9",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"b0",x"68",x"40",x"20",x"00",x"20",x"68",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"d0",x"a8",x"60",x"80",x"80",x"80",x"60",x"60",x"80",x"a0",x"a0",x"c0",x"80",x"40",x"00",x"00",x"20",x"80",x"c9",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"d6",x"b2",x"ad",x"89",x"64",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"a0",x"a4",x"c4",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"64",x"64",x"64",x"84",x"88",x"a9",x"a9",x"c9",x"c9",x"c9",x"c5",x"c5",x"c4",x"a0",x"a0",x"80",x"80",x"60",x"60",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a4",x"a8",x"ac",x"b0",x"b0",x"b0",x"b0",x"b0",x"d4",x"d8",x"f8",x"f9",x"f9",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"b0",x"88",x"44",x"20",x"00",x"20",x"48",x"6c",x"8c",x"8c",x"8c",x"b0",x"b0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d0",x"a8",x"60",x"60",x"80",x"80",x"80",x"60",x"60",x"80",x"a0",x"c0",x"a0",x"60",x"20",x"00",x"20",x"60",x"a5",x"d2",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"d2",x"ad",x"89",x"64",x"60",x"40",x"40",x"40",x"40",x"44",x"64",x"84",x"a4",x"c4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"40",x"64",x"64",x"64",x"88",x"a9",x"c9",x"e9",x"e5",x"e9",x"e9",x"e5",x"c4",x"a0",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"a0",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"c0",x"e0",x"c0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a4",x"a8",x"8c",x"b0",x"b0",x"b0",x"b0",x"b0",x"d4",x"d4",x"f8",x"f8",x"f9",x"f9",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"8c",x"44",x"20",x"00",x"20",x"44",x"68",x"8c",x"8c",x"8c",x"8c",x"b0",x"d0",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"ac",x"84",x"60",x"80",x"80",x"80",x"60",x"60",x"60",x"80",x"a0",x"c0",x"80",x"40",x"20",x"20",x"40",x"60",x"89",x"d2",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"d2",x"d2",x"ad",x"89",x"64",x"64",x"60",x"60",x"60",x"60",x"80",x"80",x"a0",x"a0",x"a4",x"c4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"64",x"64",x"64",x"84",x"a4",x"a9",x"c5",x"c5",x"c5",x"c5",x"c4",x"c4",x"c4",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"c0",x"c0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"c0",x"c0",x"a0",x"a0",x"80",x"84",x"8c",x"b0",x"b0",x"b0",x"b0",x"b0",x"d4",x"d4",x"f8",x"f8",x"f8",x"f9",x"fc",x"fc",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"ac",x"44",x"20",x"20",x"20",x"44",x"68",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"b0",x"68",x"60",x"80",x"80",x"80",x"60",x"60",x"60",x"80",x"a0",x"a0",x"a0",x"80",x"40",x"20",x"20",x"40",x"60",x"ad",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"f6",x"ce",x"a9",x"85",x"84",x"60",x"40",x"40",x"40",x"40",x"60",x"80",x"a4",x"c4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"80",x"80",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"44",x"64",x"64",x"84",x"88",x"a9",x"c9",x"e5",x"e5",x"e5",x"e4",x"c0",x"a0",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"60",x"80",x"a0",x"80",x"80",x"a0",x"c0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"a0",x"c0",x"c0",x"c0",x"a0",x"c0",x"e0",x"c0",x"a0",x"a0",x"e0",x"c0",x"a0",x"a0",x"a0",x"a0",x"c0",x"a0",x"a0",x"80",x"84",x"88",x"8c",x"b0",x"b0",x"b0",x"b0",x"b4",x"d4",x"d4",x"f8",x"f8",x"f9",x"f9",x"fc",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"b0",x"64",x"20",x"20",x"20",x"44",x"68",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"b0",x"8c",x"64",x"60",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"a0",x"a0",x"60",x"40",x"20",x"20",x"40",x"85",x"d6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"d2",x"ad",x"ad",x"a9",x"64",x"64",x"40",x"40",x"60",x"60",x"60",x"80",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"64",x"84",x"84",x"a4",x"a4",x"c4",x"c4",x"c4",x"c4",x"c4",x"a4",x"a0",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"64",x"88",x"8c",x"90",x"b0",x"b0",x"b0",x"b4",x"d4",x"d4",x"f8",x"f8",x"f8",x"f9",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"b0",x"64",x"20",x"20",x"40",x"40",x"64",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"d0",x"8c",x"84",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"80",x"40",x"00",x"00",x"40",x"60",x"89",x"d6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"d2",x"ad",x"89",x"84",x"60",x"60",x"40",x"40",x"40",x"60",x"60",x"80",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"40",x"40",x"64",x"64",x"64",x"84",x"a4",x"c4",x"c4",x"e4",x"e4",x"e0",x"c0",x"a0",x"80",x"60",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"a0",x"80",x"80",x"a0",x"c0",x"a0",x"80",x"a0",x"c0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"a0",x"c0",x"c0",x"c0",x"a0",x"a0",x"e0",x"c0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"a0",x"a0",x"a0",x"80",x"60",x"60",x"68",x"8c",x"8c",x"b0",x"b0",x"b0",x"b0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f9",x"f9",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f4",x"d0",x"68",x"40",x"40",x"40",x"40",x"44",x"88",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"ac",x"88",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"20",x"00",x"40",x"40",x"60",x"ad",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"f2",x"cd",x"a9",x"a9",x"84",x"64",x"60",x"40",x"40",x"40",x"60",x"80",x"a0",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"40",x"40",x"44",x"64",x"64",x"84",x"a4",x"c5",x"c5",x"e5",x"e4",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"a0",x"80",x"80",x"60",x"40",x"64",x"68",x"8c",x"b0",x"b0",x"b0",x"b0",x"b0",x"d4",x"d4",x"f8",x"f8",x"f9",x"f9",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"88",x"40",x"40",x"40",x"40",x"44",x"68",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d0",x"88",x"64",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"40",x"20",x"20",x"20",x"40",x"89",x"d6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"d2",x"cd",x"a9",x"a0",x"80",x"80",x"60",x"60",x"60",x"60",x"40",x"60",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"44",x"44",x"64",x"84",x"a4",x"c4",x"e5",x"e5",x"e5",x"e5",x"e0",x"c0",x"a0",x"80",x"60",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"a0",x"a0",x"c0",x"c0",x"c0",x"a0",x"c0",x"c0",x"c0",x"a0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"c0",x"c0",x"80",x"a0",x"c0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"40",x"44",x"68",x"8c",x"b0",x"b0",x"b0",x"b0",x"b0",x"d4",x"d4",x"f4",x"f8",x"f9",x"f9",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"8c",x"64",x"40",x"40",x"20",x"40",x"68",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f0",x"ac",x"64",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"40",x"20",x"20",x"20",x"64",x"ad",x"f7",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"db",x"d2",x"ad",x"a9",x"89",x"84",x"64",x"40",x"40",x"40",x"60",x"80",x"80",x"a0",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"40",x"40",x"40",x"44",x"64",x"64",x"84",x"a4",x"c5",x"c5",x"e4",x"e4",x"c4",x"c4",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"40",x"44",x"48",x"8c",x"b0",x"b0",x"b0",x"b0",x"b0",x"d4",x"d4",x"f4",x"f8",x"f9",x"f9",x"f9",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"ac",x"64",x"40",x"40",x"20",x"20",x"68",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"ac",x"a4",x"a0",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"40",x"20",x"00",x"20",x"40",x"84",x"d2",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"b2",x"b2",x"89",x"80",x"60",x"60",x"40",x"40",x"40",x"40",x"60",x"80",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"44",x"64",x"84",x"a4",x"c5",x"e5",x"e5",x"e5",x"e4",x"c0",x"a0",x"80",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"60",x"40",x"40",x"40",x"44",x"8c",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"d4",x"d4",x"f8",x"f9",x"f9",x"f9",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"ac",x"88",x"40",x"20",x"20",x"20",x"44",x"68",x"8c",x"8c",x"8c",x"ac",x"b0",x"b0",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"d8",x"d4",x"d0",x"c8",x"a0",x"80",x"80",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"20",x"20",x"20",x"20",x"40",x"a9",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"f2",x"cd",x"a9",x"84",x"64",x"44",x"40",x"40",x"40",x"60",x"60",x"80",x"80",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"64",x"64",x"84",x"a4",x"a4",x"c5",x"c5",x"e5",x"e4",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"a0",x"c0",x"c0",x"c0",x"a0",x"c0",x"c0",x"c0",x"a0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"60",x"60",x"40",x"40",x"20",x"40",x"68",x"8c",x"b0",x"b0",x"b0",x"b0",x"b0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d0",x"88",x"64",x"20",x"20",x"20",x"44",x"68",x"6c",x"8c",x"8c",x"8c",x"b0",x"b0",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"d0",x"ac",x"84",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"20",x"00",x"20",x"40",x"84",x"d2",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"d6",x"d2",x"cd",x"a9",x"80",x"60",x"60",x"40",x"40",x"40",x"60",x"60",x"80",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"60",x"60",x"40",x"40",x"40",x"44",x"44",x"64",x"84",x"84",x"a4",x"c5",x"c5",x"e5",x"e5",x"e4",x"c0",x"a0",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"00",x"20",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"68",x"8c",x"8c",x"90",x"90",x"b0",x"b0",x"d0",x"d4",x"d4",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"ac",x"64",x"20",x"20",x"40",x"44",x"68",x"68",x"8c",x"8c",x"8c",x"90",x"b0",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"b0",x"88",x"64",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"60",x"40",x"00",x"20",x"40",x"60",x"a9",x"d6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"f7",x"d2",x"cd",x"a9",x"84",x"64",x"60",x"40",x"20",x"40",x"40",x"60",x"80",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"40",x"40",x"40",x"60",x"60",x"a4",x"c4",x"c5",x"e5",x"c5",x"c4",x"c4",x"a4",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"60",x"60",x"80",x"60",x"60",x"80",x"80",x"a0",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"c0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"a0",x"a0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"a0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"c0",x"a0",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"60",x"60",x"60",x"80",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"64",x"8c",x"8c",x"90",x"b0",x"b0",x"b0",x"b0",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"ac",x"64",x"20",x"20",x"40",x"44",x"68",x"68",x"8c",x"8c",x"8c",x"90",x"b0",x"b0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"b0",x"88",x"84",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"40",x"20",x"20",x"20",x"40",x"64",x"b2",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"fb",x"d6",x"d2",x"ad",x"a9",x"80",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"80",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"60",x"60",x"60",x"80",x"a0",x"c4",x"c5",x"e5",x"c4",x"c0",x"a0",x"80",x"60",x"20",x"00",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"c0",x"a0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"64",x"68",x"8c",x"8c",x"b0",x"b0",x"b0",x"b0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"ac",x"64",x"40",x"20",x"40",x"40",x"44",x"68",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d0",x"ac",x"84",x"84",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"60",x"40",x"20",x"20",x"20",x"40",x"ad",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"f6",x"d2",x"c9",x"a5",x"a4",x"84",x"60",x"40",x"40",x"40",x"40",x"60",x"80",x"a0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"40",x"20",x"20",x"40",x"80",x"a0",x"c0",x"c0",x"e1",x"e1",x"e0",x"c0",x"a0",x"80",x"60",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"40",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"a0",x"c0",x"c0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"a0",x"c0",x"e0",x"e0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"c0",x"a0",x"80",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"a0",x"80",x"60",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"60",x"80",x"a0",x"80",x"60",x"80",x"80",x"60",x"40",x"60",x"60",x"40",x"40",x"44",x"68",x"8c",x"8c",x"b0",x"b0",x"b0",x"b0",x"b0",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d0",x"64",x"40",x"20",x"20",x"40",x"44",x"68",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"d0",x"ac",x"88",x"84",x"84",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"20",x"20",x"20",x"85",x"f2",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"fa",x"d6",x"d2",x"ad",x"a9",x"80",x"60",x"60",x"60",x"60",x"40",x"40",x"60",x"80",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"64",x"80",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"80",x"60",x"40",x"40",x"20",x"20",x"20",x"40",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"a0",x"a0",x"80",x"a0",x"c0",x"c0",x"c0",x"a0",x"a0",x"c0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"c0",x"e0",x"c0",x"c0",x"a0",x"c0",x"e0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"60",x"80",x"80",x"80",x"60",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"60",x"40",x"60",x"60",x"40",x"40",x"40",x"64",x"88",x"8c",x"b0",x"b0",x"b0",x"b0",x"b0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d0",x"88",x"40",x"40",x"20",x"20",x"44",x"68",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"b0",x"ac",x"88",x"84",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"40",x"20",x"00",x"20",x"60",x"c9",x"f6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d2",x"c9",x"a5",x"84",x"80",x"60",x"40",x"20",x"00",x"40",x"80",x"a0",x"a0",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"20",x"20",x"40",x"40",x"60",x"84",x"a4",x"c4",x"e0",x"e0",x"c0",x"c0",x"a0",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"00",x"20",x"20",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"40",x"60",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"a0",x"a0",x"a0",x"e0",x"c0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"c0",x"c0",x"80",x"80",x"c0",x"a0",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"a0",x"80",x"60",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"60",x"60",x"80",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"44",x"68",x"8c",x"ac",x"b0",x"b0",x"b0",x"b0",x"d0",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d0",x"88",x"40",x"40",x"20",x"20",x"44",x"68",x"6c",x"6c",x"8c",x"8c",x"8c",x"b0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d0",x"ac",x"88",x"84",x"84",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"20",x"00",x"20",x"40",x"80",x"d2",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"fa",x"d6",x"d2",x"ad",x"a9",x"80",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"60",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"80",x"a4",x"a4",x"c0",x"c0",x"c0",x"c0",x"a0",x"80",x"60",x"40",x"20",x"20",x"20",x"20",x"40",x"40",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"c0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"60",x"60",x"60",x"80",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"68",x"8c",x"8c",x"b0",x"b0",x"b0",x"b0",x"b0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"8c",x"64",x"40",x"20",x"20",x"40",x"68",x"68",x"6c",x"6c",x"8c",x"8c",x"b0",x"b0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d0",x"ac",x"88",x"84",x"84",x"84",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"20",x"20",x"20",x"20",x"60",x"ad",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f2",x"c9",x"a9",x"84",x"80",x"60",x"40",x"40",x"40",x"60",x"60",x"80",x"a0",x"c0",x"e0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"20",x"40",x"60",x"64",x"84",x"a4",x"c4",x"e4",x"e0",x"e0",x"c0",x"a0",x"80",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"60",x"60",x"80",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"c0",x"c0",x"a0",x"c0",x"e0",x"c0",x"c0",x"a0",x"a0",x"c0",x"c0",x"a0",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"60",x"40",x"60",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"40",x"20",x"20",x"64",x"88",x"8c",x"90",x"90",x"b0",x"b0",x"b0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"ac",x"68",x"40",x"20",x"20",x"20",x"64",x"68",x"68",x"6c",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"b0",x"88",x"84",x"84",x"84",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"40",x"20",x"20",x"20",x"40",x"89",x"d2",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"d6",x"b2",x"ad",x"89",x"84",x"60",x"60",x"40",x"60",x"60",x"60",x"80",x"80",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"a0",x"a4",x"c4",x"c4",x"c0",x"a0",x"a0",x"80",x"60",x"40",x"40",x"20",x"20",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"c0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"84",x"a4",x"a4",x"a4",x"a8",x"a8",x"a8",x"a8",x"84",x"88",x"a8",x"88",x"84",x"84",x"84",x"84",x"84",x"84",x"64",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"40",x"20",x"20",x"64",x"68",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"d0",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"b0",x"88",x"40",x"20",x"20",x"20",x"44",x"68",x"68",x"6c",x"8c",x"8c",x"8c",x"b0",x"d0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"8c",x"88",x"88",x"84",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"40",x"20",x"20",x"20",x"64",x"ad",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"f2",x"ce",x"a9",x"84",x"64",x"60",x"40",x"20",x"20",x"40",x"40",x"80",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"60",x"40",x"40",x"20",x"20",x"40",x"40",x"60",x"80",x"c0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"60",x"40",x"20",x"20",x"20",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"40",x"40",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"a0",x"c0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"a0",x"c0",x"c0",x"c0",x"a0",x"c0",x"e0",x"c0",x"a0",x"a0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"a4",x"c8",x"a8",x"a8",x"cc",x"f0",x"f0",x"f0",x"f0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f5",x"f4",x"f0",x"d0",x"d0",x"cc",x"ac",x"88",x"84",x"84",x"84",x"60",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"a0",x"80",x"40",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"44",x"48",x"88",x"8c",x"8c",x"90",x"b0",x"b0",x"b0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d0",x"8c",x"40",x"20",x"20",x"20",x"44",x"48",x"68",x"68",x"6c",x"8c",x"8c",x"b0",x"b0",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"8c",x"88",x"88",x"89",x"84",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"60",x"20",x"20",x"20",x"40",x"89",x"d6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"d6",x"b2",x"ad",x"89",x"84",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"60",x"60",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"60",x"40",x"40",x"20",x"20",x"40",x"40",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"a0",x"a0",x"a4",x"a8",x"a8",x"a8",x"cc",x"d0",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d0",x"ac",x"ac",x"ac",x"a8",x"84",x"84",x"80",x"80",x"60",x"60",x"60",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"44",x"68",x"8c",x"8c",x"8c",x"ac",x"b0",x"b0",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d0",x"ac",x"44",x"20",x"20",x"20",x"40",x"44",x"68",x"68",x"68",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d0",x"ac",x"88",x"88",x"84",x"84",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"a0",x"60",x"40",x"20",x"20",x"40",x"64",x"d2",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"ce",x"a9",x"84",x"64",x"40",x"40",x"40",x"60",x"60",x"80",x"80",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"40",x"20",x"20",x"40",x"60",x"80",x"a0",x"c0",x"e0",x"e0",x"e1",x"e0",x"a0",x"80",x"60",x"60",x"40",x"40",x"40",x"60",x"60",x"80",x"80",x"60",x"60",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"c0",x"a0",x"c0",x"e0",x"c0",x"a0",x"a0",x"c0",x"a0",x"80",x"80",x"a0",x"a4",x"a4",x"cc",x"d0",x"f4",x"f4",x"f4",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f0",x"cc",x"ac",x"88",x"64",x"60",x"60",x"60",x"40",x"60",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"20",x"20",x"40",x"64",x"68",x"6c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"ac",x"44",x"20",x"20",x"20",x"20",x"44",x"68",x"68",x"68",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"b0",x"8c",x"68",x"64",x"84",x"84",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"80",x"a0",x"80",x"40",x"20",x"20",x"20",x"40",x"ad",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"d7",x"d2",x"d2",x"ad",x"a9",x"84",x"64",x"60",x"40",x"60",x"60",x"60",x"80",x"a0",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"c0",x"a0",x"80",x"a0",x"a0",x"a0",x"a4",x"a8",x"cc",x"cc",x"d0",x"f4",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f4",x"d4",x"d0",x"ac",x"a8",x"84",x"84",x"60",x"60",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"20",x"40",x"40",x"68",x"6c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"ac",x"64",x"20",x"20",x"20",x"20",x"44",x"48",x"68",x"68",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"b0",x"8c",x"64",x"64",x"85",x"84",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"60",x"40",x"20",x"20",x"40",x"8d",x"d7",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"d6",x"b2",x"8d",x"64",x"64",x"40",x"40",x"40",x"40",x"40",x"60",x"80",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"60",x"80",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"60",x"40",x"20",x"20",x"20",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"84",x"a8",x"cc",x"f0",x"f4",x"f8",x"f9",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f4",x"d0",x"ac",x"a8",x"84",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"20",x"40",x"68",x"68",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"b0",x"64",x"20",x"20",x"20",x"20",x"44",x"48",x"68",x"68",x"68",x"8c",x"8c",x"b0",x"d0",x"d0",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"b0",x"8c",x"64",x"40",x"85",x"a5",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"40",x"20",x"20",x"20",x"69",x"d6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"f6",x"d2",x"d2",x"ad",x"89",x"69",x"64",x"40",x"40",x"40",x"60",x"60",x"80",x"a0",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"a0",x"a0",x"a0",x"a0",x"c0",x"a0",x"a0",x"a0",x"80",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a4",x"c8",x"cc",x"d0",x"f4",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f4",x"d0",x"ac",x"88",x"84",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"20",x"40",x"64",x"68",x"8c",x"8c",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"68",x"40",x"20",x"20",x"20",x"20",x"48",x"68",x"68",x"68",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"b0",x"68",x"44",x"85",x"85",x"84",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"60",x"20",x"00",x"20",x"64",x"ad",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"ce",x"c9",x"a4",x"80",x"60",x"40",x"40",x"40",x"40",x"60",x"80",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"60",x"60",x"80",x"a0",x"a0",x"c0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"40",x"40",x"20",x"20",x"20",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"a4",x"cc",x"f4",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f4",x"d0",x"a8",x"84",x"80",x"60",x"60",x"80",x"80",x"60",x"80",x"80",x"60",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"60",x"64",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"f4",x"d0",x"88",x"64",x"40",x"20",x"20",x"20",x"44",x"68",x"68",x"68",x"8c",x"8c",x"ac",x"b0",x"d0",x"d0",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"b0",x"8c",x"64",x"64",x"65",x"64",x"84",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"80",x"60",x"40",x"00",x"00",x"40",x"84",x"d6",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"f6",x"d2",x"ae",x"ad",x"89",x"84",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"a0",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"60",x"80",x"80",x"a0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"a0",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a4",x"c8",x"cc",x"f4",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f4",x"d0",x"ac",x"a8",x"84",x"80",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"64",x"68",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"d0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"f4",x"d0",x"8c",x"64",x"40",x"20",x"20",x"20",x"44",x"48",x"68",x"68",x"8c",x"8c",x"ac",x"ac",x"d0",x"d0",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"b4",x"8c",x"68",x"64",x"64",x"64",x"64",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"60",x"40",x"00",x"00",x"40",x"84",x"d2",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"ce",x"a9",x"85",x"60",x"60",x"40",x"20",x"20",x"40",x"60",x"80",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"60",x"60",x"40",x"40",x"40",x"40",x"60",x"80",x"a0",x"c0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"80",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a8",x"cc",x"f0",x"f5",x"f9",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f4",x"f4",x"d0",x"ac",x"84",x"60",x"80",x"80",x"60",x"40",x"60",x"80",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"68",x"6c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d0",x"8c",x"64",x"40",x"20",x"20",x"20",x"44",x"44",x"68",x"68",x"88",x"8c",x"8c",x"ac",x"d0",x"d0",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"8c",x"68",x"44",x"40",x"64",x"64",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"60",x"40",x"20",x"00",x"20",x"60",x"b1",x"fb",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"d2",x"d2",x"a9",x"89",x"64",x"64",x"40",x"40",x"40",x"60",x"80",x"80",x"a0",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"60",x"60",x"80",x"80",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"a4",x"c8",x"d0",x"f4",x"f9",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f4",x"f4",x"cc",x"a8",x"84",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"68",x"68",x"68",x"8c",x"8c",x"ac",x"b0",x"b0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"ac",x"68",x"40",x"20",x"20",x"20",x"44",x"44",x"68",x"68",x"68",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"b0",x"8c",x"44",x"20",x"44",x"64",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"60",x"40",x"20",x"00",x"20",x"40",x"89",x"d6",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"d2",x"ad",x"a5",x"80",x"60",x"40",x"40",x"40",x"40",x"40",x"80",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"20",x"24",x"60",x"80",x"a0",x"c0",x"e0",x"e0",x"e0",x"c0",x"a0",x"60",x"40",x"40",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"a0",x"c0",x"a0",x"80",x"a0",x"c0",x"c0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"c0",x"a0",x"c0",x"c0",x"a0",x"a0",x"a0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"60",x"80",x"80",x"60",x"84",x"ac",x"f4",x"f4",x"f8",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f4",x"f0",x"88",x"40",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"20",x"40",x"44",x"68",x"68",x"8c",x"8c",x"8c",x"ac",x"b0",x"b0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"ac",x"88",x"40",x"20",x"20",x"20",x"20",x"44",x"48",x"68",x"68",x"88",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"b0",x"8c",x"44",x"20",x"24",x"44",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"20",x"20",x"20",x"40",x"85",x"b2",x"fb",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"d2",x"ad",x"a9",x"89",x"84",x"64",x"60",x"40",x"60",x"60",x"80",x"80",x"a0",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"80",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"88",x"ac",x"f4",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"d0",x"ac",x"84",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"60",x"40",x"40",x"40",x"44",x"64",x"68",x"8c",x"8c",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"88",x"40",x"20",x"20",x"20",x"20",x"44",x"44",x"68",x"68",x"68",x"88",x"8c",x"b0",x"d0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"8c",x"44",x"20",x"24",x"44",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"40",x"20",x"20",x"20",x"60",x"a9",x"fb",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"f6",x"d2",x"cd",x"a9",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"80",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"60",x"60",x"80",x"a0",x"c0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"40",x"20",x"20",x"20",x"20",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"40",x"40",x"40",x"20",x"20",x"20",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"60",x"60",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"a0",x"a0",x"c0",x"c0",x"c0",x"a0",x"c0",x"e0",x"c0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"60",x"64",x"d0",x"f4",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f4",x"ac",x"64",x"60",x"80",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"44",x"68",x"8c",x"8c",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d0",x"8c",x"44",x"20",x"20",x"20",x"20",x"44",x"44",x"68",x"68",x"68",x"88",x"8c",x"ac",x"d0",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"b0",x"48",x"24",x"24",x"20",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"40",x"20",x"20",x"20",x"40",x"85",x"d6",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"d2",x"cd",x"a9",x"89",x"64",x"64",x"40",x"40",x"60",x"60",x"80",x"a0",x"a0",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"80",x"84",x"84",x"80",x"60",x"40",x"40",x"40",x"20",x"40",x"60",x"80",x"80",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"88",x"d0",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"d4",x"ac",x"84",x"80",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"44",x"68",x"88",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d0",x"ac",x"64",x"20",x"20",x"20",x"20",x"44",x"44",x"68",x"68",x"68",x"68",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"b0",x"6c",x"44",x"04",x"20",x"40",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"20",x"00",x"40",x"84",x"d6",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"db",x"da",x"d2",x"c9",x"a5",x"80",x"60",x"40",x"40",x"40",x"40",x"40",x"60",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"84",x"84",x"88",x"a8",x"88",x"88",x"64",x"40",x"44",x"24",x"20",x"40",x"80",x"c0",x"c0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"40",x"20",x"20",x"20",x"40",x"40",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"c0",x"a0",x"c0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"c0",x"c0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"84",x"88",x"d0",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"ac",x"84",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"44",x"68",x"68",x"8c",x"8c",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"ac",x"64",x"40",x"20",x"20",x"20",x"20",x"44",x"68",x"68",x"68",x"68",x"8c",x"ac",x"b0",x"d0",x"d0",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"b0",x"8c",x"48",x"04",x"00",x"40",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"40",x"20",x"00",x"20",x"60",x"d2",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"f2",x"cd",x"a9",x"89",x"64",x"60",x"40",x"40",x"40",x"60",x"80",x"80",x"a0",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a8",x"ac",x"d0",x"d4",x"d4",x"d4",x"f4",x"d4",x"d4",x"d0",x"cc",x"ac",x"a8",x"80",x"a0",x"c0",x"c0",x"c0",x"a0",x"80",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"c0",x"c0",x"c0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"c0",x"c0",x"a0",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"80",x"80",x"80",x"80",x"80",x"84",x"ac",x"d4",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"cc",x"84",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"64",x"68",x"88",x"8c",x"8c",x"8c",x"8c",x"b0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"b0",x"68",x"40",x"20",x"20",x"20",x"20",x"44",x"44",x"68",x"68",x"68",x"8c",x"8c",x"b0",x"b0",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"6c",x"24",x"00",x"20",x"40",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"20",x"00",x"20",x"60",x"d2",x"fb",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"d2",x"cd",x"a9",x"84",x"60",x"60",x"40",x"40",x"40",x"40",x"60",x"80",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"a0",x"a8",x"d0",x"f4",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f1",x"ec",x"e8",x"c0",x"c0",x"a0",x"a0",x"80",x"40",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"c0",x"a0",x"c0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"80",x"80",x"c0",x"c0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"a0",x"80",x"60",x"80",x"80",x"80",x"88",x"d4",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f8",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"a8",x"80",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"64",x"68",x"68",x"88",x"8c",x"8c",x"8c",x"b0",x"b0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"b0",x"88",x"44",x"20",x"20",x"20",x"20",x"44",x"44",x"68",x"68",x"68",x"88",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"8c",x"24",x"00",x"20",x"40",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"20",x"00",x"20",x"60",x"ad",x"fb",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"f2",x"cd",x"c9",x"a4",x"84",x"60",x"40",x"40",x"40",x"40",x"60",x"80",x"a0",x"a0",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"a8",x"cc",x"f4",x"f9",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f4",x"d0",x"a8",x"60",x"40",x"60",x"60",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"a8",x"d0",x"f4",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"f4",x"f4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d0",x"ac",x"84",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"64",x"68",x"68",x"8c",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"88",x"64",x"20",x"20",x"20",x"20",x"44",x"44",x"68",x"68",x"68",x"68",x"8c",x"8c",x"b0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"90",x"48",x"20",x"24",x"44",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"20",x"00",x"20",x"40",x"a9",x"f6",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"db",x"d6",x"d2",x"cd",x"c5",x"a0",x"80",x"60",x"40",x"40",x"40",x"40",x"60",x"60",x"80",x"c4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"88",x"d0",x"f4",x"f9",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"d8",x"b0",x"48",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"c0",x"e0",x"c0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"a0",x"80",x"80",x"80",x"a0",x"a0",x"80",x"60",x"80",x"80",x"60",x"88",x"d0",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"f5",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"d0",x"d0",x"d0",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d0",x"a8",x"84",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"64",x"68",x"68",x"88",x"8c",x"8c",x"8c",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"8c",x"64",x"20",x"20",x"20",x"20",x"44",x"44",x"48",x"68",x"68",x"68",x"88",x"8c",x"ac",x"b0",x"d0",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"b0",x"68",x"24",x"24",x"24",x"64",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"20",x"00",x"00",x"40",x"a9",x"f2",x"fb",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d7",x"d6",x"ae",x"a9",x"84",x"64",x"60",x"40",x"40",x"40",x"60",x"60",x"80",x"a0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"40",x"20",x"44",x"b0",x"d8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"d4",x"b0",x"88",x"40",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"a8",x"d0",x"f4",x"f8",x"fc",x"fc",x"fc",x"fc",x"f9",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f4",x"d4",x"d4",x"d4",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"ac",x"b0",x"b0",x"b0",x"b0",x"b0",x"d0",x"d0",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d0",x"88",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"44",x"64",x"68",x"68",x"8c",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"8c",x"64",x"20",x"20",x"20",x"20",x"40",x"44",x"44",x"68",x"68",x"68",x"68",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"b0",x"68",x"44",x"24",x"24",x"64",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"20",x"00",x"00",x"40",x"85",x"ce",x"fb",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"d6",x"b2",x"8e",x"89",x"64",x"60",x"60",x"40",x"40",x"40",x"40",x"60",x"80",x"a4",x"c4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"20",x"68",x"d4",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f4",x"b0",x"64",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"88",x"d0",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"f9",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f5",x"d4",x"d4",x"b0",x"b0",x"b0",x"90",x"90",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"ac",x"b0",x"b0",x"b0",x"b0",x"b0",x"d0",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"ac",x"88",x"60",x"40",x"40",x"40",x"40",x"40",x"44",x"64",x"68",x"68",x"8c",x"8c",x"8c",x"ac",x"b0",x"d0",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"ac",x"68",x"40",x"20",x"20",x"20",x"40",x"44",x"44",x"48",x"68",x"68",x"68",x"8c",x"8c",x"b0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"b0",x"8c",x"68",x"24",x"24",x"64",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"40",x"00",x"00",x"20",x"84",x"c9",x"fb",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"f2",x"cd",x"c9",x"a4",x"64",x"40",x"20",x"20",x"40",x"60",x"60",x"84",x"a4",x"c4",x"c4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"60",x"40",x"20",x"20",x"20",x"40",x"60",x"80",x"a8",x"d0",x"f8",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fd",x"fd",x"fe",x"fe",x"fe",x"fd",x"fd",x"f8",x"f8",x"f8",x"d4",x"ac",x"88",x"40",x"20",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a4",x"cc",x"f4",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"f9",x"f9",x"f5",x"d5",x"d4",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"6c",x"6c",x"6c",x"6c",x"68",x"68",x"68",x"68",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"ac",x"ac",x"ac",x"b0",x"b0",x"d0",x"d4",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"cc",x"88",x"60",x"40",x"40",x"40",x"40",x"40",x"44",x"64",x"68",x"6c",x"8c",x"8c",x"8c",x"ac",x"d0",x"d0",x"d0",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"d0",x"8c",x"44",x"20",x"20",x"20",x"40",x"44",x"44",x"44",x"44",x"68",x"68",x"88",x"8c",x"b0",x"d0",x"d0",x"d0",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"ac",x"88",x"24",x"24",x"84",x"a4",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"60",x"20",x"20",x"20",x"40",x"85",x"f6",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"d6",x"d2",x"ad",x"a9",x"84",x"80",x"60",x"60",x"40",x"40",x"40",x"60",x"84",x"a4",x"c4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"60",x"80",x"a4",x"ec",x"f4",x"f8",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fd",x"fd",x"fe",x"fe",x"ff",x"fe",x"fd",x"f8",x"f8",x"f8",x"f4",x"d0",x"88",x"40",x"20",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"ac",x"f0",x"f8",x"fc",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f9",x"d4",x"d4",x"d0",x"b0",x"8c",x"8c",x"8c",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"68",x"68",x"68",x"68",x"68",x"6c",x"6c",x"6c",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"ac",x"b0",x"b0",x"d0",x"d4",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d0",x"ac",x"64",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"68",x"6c",x"6c",x"8c",x"8c",x"ac",x"b0",x"d0",x"d0",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"d0",x"ac",x"64",x"40",x"40",x"20",x"40",x"40",x"44",x"44",x"44",x"48",x"68",x"88",x"8c",x"b0",x"d0",x"d0",x"d0",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"d0",x"8c",x"24",x"24",x"84",x"a4",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"60",x"40",x"20",x"20",x"40",x"60",x"d6",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"da",x"d2",x"cd",x"a9",x"a4",x"80",x"60",x"40",x"20",x"40",x"44",x"64",x"a4",x"c4",x"c4",x"e5",x"e5",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"40",x"20",x"40",x"60",x"80",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"c4",x"f0",x"f4",x"f8",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fd",x"fd",x"fe",x"fe",x"fd",x"f9",x"f8",x"f8",x"f8",x"f4",x"d0",x"8c",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"a0",x"a0",x"60",x"80",x"a0",x"c0",x"80",x"60",x"80",x"a0",x"80",x"80",x"80",x"80",x"a0",x"80",x"80",x"80",x"a8",x"d0",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"d5",x"d4",x"b0",x"b0",x"8c",x"8c",x"8c",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"48",x"48",x"68",x"68",x"68",x"68",x"68",x"6c",x"6c",x"6c",x"6c",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"ac",x"b0",x"b0",x"b0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"ac",x"84",x"60",x"40",x"40",x"40",x"40",x"40",x"44",x"68",x"68",x"68",x"68",x"8c",x"ac",x"b0",x"d0",x"d0",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"d0",x"ac",x"64",x"40",x"20",x"20",x"20",x"40",x"44",x"44",x"44",x"48",x"68",x"68",x"8c",x"b0",x"d0",x"d0",x"d0",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"d0",x"8c",x"48",x"44",x"84",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"60",x"40",x"20",x"20",x"40",x"84",x"d6",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"d6",x"b2",x"8d",x"89",x"84",x"80",x"60",x"60",x"60",x"40",x"40",x"64",x"84",x"a4",x"c4",x"e4",x"e5",x"e5",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"60",x"40",x"40",x"60",x"80",x"a0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a4",x"f0",x"f8",x"f8",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"f9",x"f8",x"f8",x"f4",x"d4",x"d4",x"8c",x"44",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"40",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a4",x"cc",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"d4",x"d4",x"b0",x"8c",x"8c",x"8c",x"68",x"68",x"68",x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"6c",x"8c",x"8c",x"8c",x"ac",x"ac",x"b0",x"b0",x"b0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d0",x"a8",x"64",x"40",x"40",x"40",x"40",x"40",x"44",x"68",x"68",x"68",x"68",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"d0",x"ac",x"64",x"40",x"20",x"20",x"20",x"40",x"44",x"44",x"44",x"48",x"68",x"68",x"8c",x"ac",x"d0",x"d0",x"d0",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"d0",x"ac",x"48",x"44",x"64",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"60",x"40",x"20",x"20",x"40",x"84",x"d6",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f2",x"cd",x"c9",x"a5",x"60",x"40",x"40",x"40",x"40",x"40",x"64",x"84",x"a4",x"c4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"60",x"60",x"40",x"20",x"20",x"20",x"20",x"60",x"80",x"a0",x"a0",x"e0",x"e0",x"e0",x"e0",x"a0",x"80",x"60",x"40",x"40",x"68",x"d4",x"f8",x"f8",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"f9",x"f9",x"f8",x"f8",x"f4",x"d4",x"d4",x"b0",x"44",x"20",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"c0",x"c0",x"a0",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"c0",x"a0",x"80",x"80",x"80",x"a0",x"c0",x"80",x"80",x"80",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"60",x"80",x"a0",x"a0",x"80",x"80",x"84",x"cc",x"f0",x"f5",x"f9",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"d4",x"b0",x"b0",x"8c",x"8c",x"6c",x"6c",x"68",x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"68",x"68",x"8c",x"8c",x"8c",x"8c",x"8c",x"ac",x"b0",x"b0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d0",x"88",x"60",x"40",x"40",x"40",x"40",x"44",x"68",x"68",x"68",x"68",x"68",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d0",x"d0",x"ac",x"68",x"40",x"20",x"20",x"20",x"20",x"44",x"44",x"44",x"48",x"68",x"68",x"8c",x"ac",x"b0",x"d0",x"d0",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"d0",x"ac",x"6c",x"48",x"64",x"80",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"60",x"40",x"20",x"20",x"40",x"84",x"d2",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"d6",x"d6",x"d2",x"ad",x"a9",x"84",x"80",x"60",x"60",x"60",x"60",x"60",x"64",x"84",x"a4",x"c4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"a0",x"80",x"60",x"40",x"40",x"40",x"68",x"d4",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"f9",x"f9",x"f8",x"f8",x"f4",x"d4",x"d4",x"b0",x"68",x"24",x"20",x"00",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"a0",x"80",x"80",x"80",x"a8",x"d0",x"f4",x"f9",x"f9",x"f8",x"f8",x"fc",x"fc",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"d4",x"b0",x"b0",x"8c",x"8c",x"6c",x"6c",x"68",x"68",x"48",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"48",x"48",x"68",x"68",x"68",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d0",x"ac",x"64",x"40",x"40",x"40",x"40",x"44",x"44",x"68",x"68",x"68",x"68",x"8c",x"8c",x"b0",x"d0",x"d0",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"ac",x"88",x"44",x"20",x"20",x"20",x"20",x"44",x"44",x"44",x"48",x"68",x"68",x"8c",x"ac",x"b0",x"d0",x"d0",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"8c",x"68",x"44",x"80",x"c0",x"c0",x"a0",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"40",x"20",x"20",x"40",x"60",x"d2",x"fb"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"f2",x"cd",x"a9",x"84",x"80",x"60",x"40",x"40",x"40",x"40",x"84",x"a4",x"c4",x"c4",x"c4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"80",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"20",x"20",x"20",x"40",x"60",x"80",x"a0",x"c0",x"e0",x"e0",x"c0",x"a0",x"a0",x"80",x"60",x"40",x"20",x"20",x"40",x"40",x"60",x"60",x"60",x"a8",x"f4",x"f8",x"f8",x"f8",x"f9",x"f9",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f8",x"d4",x"8c",x"44",x"20",x"20",x"20",x"20",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"c4",x"c4",x"c4",x"c4",x"e4",x"e4",x"e4",x"e4",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"c0",x"c0",x"a0",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"60",x"a0",x"c0",x"a0",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"c0",x"a0",x"60",x"80",x"a0",x"a4",x"cc",x"f4",x"f8",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f5",x"d4",x"b0",x"b0",x"8c",x"8c",x"6c",x"68",x"68",x"68",x"48",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"40",x"40",x"20",x"20",x"40",x"40",x"44",x"44",x"44",x"44",x"44",x"44",x"48",x"68",x"68",x"68",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d0",x"88",x"60",x"40",x"40",x"40",x"40",x"44",x"44",x"68",x"68",x"68",x"88",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"88",x"64",x"20",x"20",x"20",x"20",x"40",x"44",x"44",x"48",x"68",x"68",x"88",x"8c",x"ac",x"d0",x"d0",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"d0",x"ac",x"6c",x"44",x"60",x"c0",x"e0",x"c0",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"20",x"00",x"20",x"60",x"d2",x"fb"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"d6",x"d2",x"ad",x"89",x"84",x"60",x"60",x"60",x"60",x"60",x"60",x"84",x"84",x"c4",x"e4",x"e4",x"e4",x"e5",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"60",x"60",x"80",x"80",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"80",x"60",x"60",x"40",x"40",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"88",x"d4",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"8c",x"68",x"20",x"20",x"40",x"40",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c4",x"c4",x"c4",x"c8",x"c8",x"c8",x"c8",x"ec",x"ec",x"ec",x"ec",x"f0",x"f0",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"c8",x"c4",x"c4",x"c4",x"c4",x"c4",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a8",x"d0",x"f4",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"d4",x"b0",x"b0",x"8c",x"8c",x"8c",x"68",x"68",x"68",x"44",x"44",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"44",x"44",x"44",x"48",x"48",x"68",x"68",x"68",x"88",x"88",x"8c",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d0",x"ac",x"84",x"40",x"40",x"20",x"40",x"44",x"44",x"68",x"68",x"68",x"68",x"88",x"ac",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"8c",x"64",x"20",x"20",x"20",x"20",x"20",x"44",x"44",x"48",x"68",x"68",x"68",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"8c",x"48",x"64",x"c0",x"e0",x"c0",x"a0",x"60",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"20",x"00",x"20",x"60",x"d2",x"fb"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"f6",x"ee",x"c9",x"a5",x"84",x"40",x"40",x"20",x"40",x"44",x"64",x"84",x"a4",x"c5",x"e9",x"e5",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"40",x"20",x"20",x"40",x"60",x"80",x"a0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"60",x"60",x"40",x"40",x"40",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"68",x"d4",x"f8",x"d4",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"b0",x"88",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e4",x"e4",x"e8",x"ec",x"f0",x"f0",x"f4",x"f5",x"f9",x"f9",x"f9",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"cc",x"c8",x"a4",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"c0",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"a0",x"c0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"a0",x"c0",x"a0",x"80",x"80",x"a0",x"a0",x"84",x"ac",x"f4",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"d4",x"b0",x"b0",x"8c",x"8c",x"88",x"68",x"68",x"44",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"44",x"44",x"48",x"48",x"48",x"68",x"68",x"68",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"cc",x"88",x"40",x"40",x"20",x"40",x"44",x"44",x"68",x"68",x"68",x"68",x"88",x"8c",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"ac",x"68",x"40",x"20",x"20",x"20",x"20",x"44",x"44",x"48",x"68",x"68",x"68",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"8c",x"48",x"64",x"c0",x"e0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"20",x"00",x"20",x"60",x"d2",x"f6"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"d2",x"ce",x"cd",x"a9",x"84",x"84",x"64",x"60",x"60",x"60",x"64",x"84",x"84",x"a4",x"c9",x"e5",x"e5",x"e5",x"e5",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"60",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"64",x"d0",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"d0",x"ac",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c4",x"e4",x"e8",x"e8",x"ec",x"f0",x"f0",x"f4",x"f4",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f0",x"cc",x"cc",x"c8",x"a8",x"a4",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a4",x"a4",x"cc",x"f4",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"b0",x"8c",x"8c",x"68",x"68",x"68",x"64",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"44",x"44",x"44",x"48",x"68",x"68",x"68",x"68",x"8c",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d0",x"ac",x"64",x"40",x"20",x"20",x"40",x"44",x"68",x"68",x"68",x"68",x"68",x"8c",x"ac",x"b0",x"d0",x"d0",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"88",x"40",x"20",x"20",x"20",x"20",x"44",x"44",x"48",x"68",x"68",x"68",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"68",x"84",x"c0",x"e0",x"e0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"20",x"00",x"20",x"40",x"ad",x"f6"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"d2",x"ad",x"85",x"80",x"60",x"60",x"24",x"24",x"64",x"84",x"a8",x"c9",x"e9",x"e5",x"e5",x"e5",x"e5",x"e5",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"40",x"20",x"20",x"20",x"40",x"60",x"80",x"a0",x"c0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"60",x"40",x"20",x"20",x"20",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"64",x"cc",x"f4",x"d8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"d4",x"d4",x"ac",x"84",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c4",x"c4",x"c8",x"f0",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"cc",x"cc",x"a8",x"84",x"80",x"a0",x"c0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"a0",x"c0",x"a0",x"80",x"a0",x"a0",x"a0",x"80",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"c0",x"a0",x"80",x"84",x"a8",x"d0",x"f4",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"f8",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"88",x"68",x"68",x"44",x"44",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"44",x"44",x"44",x"68",x"68",x"68",x"8c",x"8c",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"ac",x"88",x"40",x"40",x"20",x"40",x"44",x"64",x"68",x"68",x"68",x"68",x"8c",x"ac",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"8c",x"44",x"20",x"20",x"20",x"20",x"20",x"44",x"44",x"68",x"68",x"68",x"88",x"8c",x"b0",x"d0",x"d0",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"b0",x"6c",x"88",x"c4",x"e0",x"e0",x"c0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"20",x"00",x"00",x"40",x"ad",x"f6"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"d2",x"d2",x"ad",x"a9",x"84",x"84",x"64",x"60",x"60",x"64",x"64",x"68",x"88",x"a9",x"c9",x"e9",x"e5",x"e5",x"e5",x"e5",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"80",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"40",x"20",x"20",x"44",x"ac",x"d4",x"d8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"d4",x"f4",x"cc",x"84",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c4",x"e8",x"ec",x"f0",x"f4",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f4",x"f4",x"f0",x"cc",x"a8",x"c4",x"a4",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"84",x"a8",x"ac",x"d0",x"f4",x"f8",x"f8",x"f9",x"fd",x"fd",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"68",x"68",x"44",x"44",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"44",x"44",x"68",x"68",x"68",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d0",x"88",x"64",x"40",x"20",x"40",x"44",x"64",x"64",x"68",x"68",x"68",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"8c",x"64",x"20",x"20",x"20",x"20",x"20",x"44",x"44",x"68",x"68",x"68",x"88",x"8c",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"b0",x"8c",x"88",x"c4",x"e0",x"e0",x"c0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"20",x"00",x"00",x"40",x"ad",x"f2"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"d2",x"a9",x"a5",x"80",x"80",x"60",x"60",x"60",x"64",x"88",x"89",x"8d",x"cd",x"e9",x"e9",x"e9",x"e9",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"40",x"40",x"40",x"40",x"60",x"80",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"40",x"20",x"20",x"44",x"8c",x"b0",x"d8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"d4",x"f4",x"d0",x"a8",x"a4",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c4",x"c8",x"ec",x"f0",x"f4",x"f9",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"fc",x"f8",x"f8",x"f5",x"f0",x"cc",x"a8",x"a4",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"80",x"a0",x"c0",x"a0",x"80",x"a0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"60",x"80",x"c0",x"c0",x"80",x"80",x"a4",x"c8",x"b0",x"d4",x"f4",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"d4",x"b0",x"b0",x"8c",x"8c",x"88",x"68",x"64",x"44",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"44",x"48",x"68",x"68",x"68",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d0",x"ac",x"64",x"40",x"20",x"20",x"40",x"44",x"44",x"64",x"68",x"68",x"68",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"ac",x"64",x"40",x"20",x"20",x"20",x"20",x"44",x"44",x"68",x"68",x"68",x"88",x"8c",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"b0",x"b0",x"ac",x"c4",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"20",x"00",x"20",x"40",x"ad",x"d2"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"db",x"d7",x"d2",x"ad",x"a9",x"a9",x"84",x"64",x"60",x"60",x"60",x"84",x"84",x"a4",x"a9",x"a9",x"c9",x"c9",x"e9",x"e9",x"e9",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"20",x"20",x"00",x"20",x"68",x"90",x"d8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f9",x"f9",x"f9",x"f8",x"d4",x"d4",x"f4",x"d0",x"c8",x"a4",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c4",x"e8",x"ec",x"f0",x"f4",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f4",x"d0",x"cc",x"c8",x"a4",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a4",x"ac",x"d0",x"d4",x"f4",x"f8",x"f9",x"fd",x"fd",x"fd",x"fd",x"fc",x"f8",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"88",x"68",x"64",x"44",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"44",x"44",x"48",x"68",x"68",x"68",x"8c",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d0",x"ac",x"88",x"40",x"20",x"20",x"20",x"44",x"44",x"44",x"68",x"68",x"68",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"ac",x"64",x"40",x"20",x"20",x"20",x"20",x"44",x"44",x"68",x"68",x"68",x"88",x"8c",x"b0",x"b0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"b0",x"b0",x"ac",x"c4",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"20",x"00",x"20",x"40",x"a9",x"d2"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"b2",x"8d",x"85",x"80",x"60",x"60",x"60",x"60",x"64",x"68",x"89",x"ad",x"cd",x"cd",x"ed",x"e9",x"e9",x"e5",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"20",x"20",x"44",x"64",x"84",x"a0",x"c0",x"e0",x"e0",x"c0",x"c0",x"a0",x"60",x"40",x"20",x"20",x"20",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"20",x"20",x"20",x"40",x"40",x"20",x"20",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"44",x"8c",x"d4",x"f8",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"fd",x"fd",x"f9",x"f8",x"d4",x"d4",x"f4",x"f0",x"cc",x"c4",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c4",x"e8",x"ec",x"f4",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"f9",x"f4",x"f0",x"cc",x"a4",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"84",x"ac",x"d4",x"f4",x"f4",x"f8",x"f9",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"b0",x"b0",x"8c",x"8c",x"68",x"64",x"44",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"24",x"44",x"44",x"68",x"68",x"68",x"88",x"8c",x"8c",x"8c",x"ac",x"b0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"d0",x"88",x"64",x"20",x"20",x"20",x"40",x"44",x"44",x"68",x"68",x"68",x"88",x"ac",x"b0",x"d0",x"d0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"b0",x"68",x"40",x"20",x"20",x"20",x"20",x"44",x"44",x"68",x"68",x"68",x"68",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"d0",x"cc",x"c8",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"60",x"80",x"80",x"80",x"a0",x"80",x"20",x"00",x"20",x"40",x"a9",x"ce"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"d2",x"ad",x"89",x"89",x"65",x"64",x"64",x"64",x"64",x"84",x"84",x"89",x"a9",x"ad",x"cd",x"cd",x"ed",x"e9",x"e9",x"e5",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"60",x"60",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"68",x"d4",x"f8",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f9",x"f8",x"f8",x"d8",x"d8",x"d4",x"d0",x"c8",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e8",x"ec",x"f0",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f4",x"f4",x"d0",x"cc",x"a4",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"84",x"a8",x"b0",x"d4",x"f4",x"f4",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f8",x"d4",x"d4",x"d0",x"b0",x"ac",x"8c",x"88",x"64",x"64",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"44",x"44",x"68",x"68",x"68",x"88",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"ac",x"64",x"40",x"20",x"20",x"20",x"44",x"44",x"64",x"68",x"68",x"68",x"8c",x"ac",x"ac",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"88",x"64",x"20",x"20",x"20",x"20",x"44",x"44",x"68",x"68",x"68",x"68",x"8c",x"8c",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"cc",x"a8",x"c4",x"e0",x"e0",x"a0",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"20",x"00",x"20",x"60",x"a9",x"d2"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"f2",x"c9",x"84",x"60",x"60",x"40",x"40",x"40",x"64",x"69",x"89",x"ad",x"cd",x"cd",x"ed",x"ed",x"ed",x"e9",x"e8",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"60",x"60",x"40",x"40",x"20",x"20",x"40",x"40",x"60",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"60",x"40",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"20",x"20",x"20",x"68",x"b4",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"d8",x"d8",x"d4",x"f0",x"e8",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e8",x"f0",x"f4",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"ff",x"ff",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"d4",x"cc",x"a4",x"a0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"c0",x"80",x"80",x"a0",x"a0",x"80",x"a0",x"c0",x"a0",x"80",x"84",x"ac",x"d0",x"d4",x"d4",x"f4",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f4",x"d0",x"d0",x"b0",x"b0",x"8c",x"8c",x"68",x"64",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"64",x"68",x"68",x"68",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"ac",x"88",x"64",x"40",x"20",x"20",x"40",x"44",x"44",x"44",x"68",x"68",x"88",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"ac",x"68",x"20",x"20",x"20",x"20",x"20",x"44",x"68",x"68",x"68",x"68",x"88",x"8c",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"d0",x"8c",x"a8",x"e0",x"e0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"20",x"00",x"20",x"60",x"ad",x"d2"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"d2",x"ad",x"a9",x"85",x"84",x"64",x"64",x"64",x"64",x"84",x"89",x"a9",x"a9",x"cd",x"cd",x"cd",x"ed",x"e9",x"e9",x"e9",x"e5",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"64",x"64",x"84",x"a4",x"c4",x"c0",x"c0",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"60",x"60",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"20",x"20",x"64",x"b0",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"d8",x"d4",x"d4",x"d0",x"cc",x"c4",x"c0",x"e0",x"e0",x"e4",x"e8",x"ec",x"f0",x"f4",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f4",x"f0",x"cc",x"c8",x"a4",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"84",x"88",x"ac",x"d0",x"d4",x"d4",x"f8",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f5",x"f9",x"f4",x"d0",x"b0",x"b0",x"b0",x"8c",x"88",x"68",x"64",x"40",x"40",x"40",x"60",x"60",x"60",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"44",x"68",x"68",x"68",x"8c",x"8c",x"8c",x"ac",x"d0",x"d0",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"b0",x"88",x"64",x"40",x"20",x"20",x"40",x"44",x"44",x"44",x"68",x"68",x"88",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"ac",x"68",x"20",x"20",x"20",x"20",x"20",x"44",x"68",x"68",x"68",x"68",x"68",x"8c",x"b0",x"b0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"f0",x"d0",x"8c",x"a8",x"e0",x"e0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"20",x"00",x"20",x"60",x"ad",x"d2"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"d6",x"d2",x"ad",x"85",x"60",x"40",x"40",x"40",x"44",x"68",x"6d",x"8d",x"ad",x"cd",x"ed",x"ed",x"ed",x"ed",x"e9",x"e9",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"40",x"40",x"60",x"60",x"84",x"a4",x"c4",x"e5",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"64",x"b0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"d4",x"d0",x"cc",x"c4",x"c0",x"e0",x"e4",x"e8",x"ec",x"f0",x"f5",x"f9",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fc",x"f8",x"f8",x"f4",x"f4",x"f4",x"d0",x"c8",x"a4",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"84",x"a8",x"ac",x"d0",x"d4",x"f4",x"f8",x"f9",x"fd",x"fd",x"fd",x"fd",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f9",x"f4",x"d0",x"b0",x"b0",x"b0",x"8c",x"88",x"64",x"64",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"60",x"60",x"60",x"40",x"60",x"60",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"44",x"64",x"68",x"68",x"88",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d0",x"b0",x"8c",x"64",x"40",x"20",x"20",x"40",x"44",x"44",x"68",x"68",x"68",x"88",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"b0",x"68",x"40",x"20",x"20",x"20",x"20",x"44",x"68",x"68",x"68",x"68",x"68",x"8c",x"b0",x"b0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"f4",x"d0",x"ac",x"a8",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"20",x"00",x"20",x"60",x"ad",x"d2"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"d2",x"c9",x"a9",x"85",x"84",x"64",x"64",x"64",x"64",x"68",x"89",x"8d",x"ad",x"d1",x"d1",x"ed",x"ed",x"ed",x"e9",x"e9",x"e9",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"40",x"40",x"40",x"64",x"84",x"a4",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"40",x"40",x"40",x"64",x"8c",x"d0",x"f4",x"f8",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f9",x"f9",x"f8",x"d4",x"d4",x"d0",x"cc",x"c8",x"e4",x"e4",x"ec",x"f0",x"f4",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fc",x"fc",x"f8",x"f8",x"f8",x"f4",x"d0",x"ac",x"a4",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"84",x"a8",x"d0",x"d0",x"d4",x"f4",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d0",x"b0",x"b0",x"ac",x"8c",x"68",x"64",x"44",x"40",x"40",x"40",x"60",x"60",x"60",x"40",x"60",x"60",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"64",x"68",x"68",x"68",x"88",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d0",x"d0",x"ac",x"64",x"40",x"20",x"20",x"40",x"44",x"44",x"68",x"68",x"68",x"88",x"8c",x"8c",x"ac",x"d0",x"d0",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"b0",x"88",x"40",x"20",x"20",x"20",x"20",x"44",x"68",x"68",x"68",x"68",x"68",x"8c",x"ac",x"b0",x"d0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"b0",x"a8",x"e4",x"e0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"60",x"80",x"60",x"20",x"00",x"20",x"60",x"ad",x"d2"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"d2",x"ad",x"a5",x"a0",x"80",x"60",x"60",x"60",x"64",x"69",x"8d",x"ad",x"d1",x"f2",x"f2",x"f2",x"ed",x"ed",x"e9",x"e9",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"40",x"40",x"40",x"44",x"84",x"a4",x"c4",x"e5",x"e1",x"e0",x"e0",x"c0",x"80",x"60",x"40",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"60",x"88",x"b0",x"f4",x"f8",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f9",x"f9",x"f8",x"d4",x"d4",x"d4",x"d0",x"cc",x"e8",x"ec",x"f0",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f8",x"d8",x"d0",x"cc",x"c4",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"80",x"80",x"c0",x"c0",x"a0",x"80",x"a0",x"a0",x"84",x"a8",x"d0",x"d4",x"d4",x"f4",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"8c",x"8c",x"68",x"64",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"60",x"80",x"40",x"40",x"60",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"60",x"60",x"60",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"44",x"64",x"68",x"68",x"88",x"8c",x"8c",x"ac",x"d0",x"d0",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d0",x"d0",x"ac",x"88",x"40",x"20",x"20",x"20",x"40",x"44",x"68",x"68",x"68",x"68",x"88",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"b0",x"8c",x"44",x"20",x"20",x"20",x"20",x"44",x"68",x"68",x"68",x"68",x"68",x"8c",x"ac",x"b0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f9",x"f8",x"f4",x"f4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"b0",x"ac",x"c8",x"e0",x"e0",x"a0",x"80",x"80",x"80",x"80",x"60",x"80",x"60",x"20",x"00",x"20",x"60",x"ad",x"d2"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"d2",x"cd",x"a9",x"85",x"84",x"64",x"64",x"69",x"69",x"89",x"8d",x"ad",x"ad",x"d1",x"d1",x"f1",x"ed",x"ed",x"ed",x"e9",x"e9",x"e5",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"60",x"64",x"84",x"a4",x"c4",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"84",x"ac",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"d4",x"d4",x"d4",x"d0",x"d0",x"f0",x"f0",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d0",x"cc",x"a4",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a8",x"ac",x"b0",x"d4",x"d4",x"f4",x"f8",x"fd",x"fd",x"fd",x"fd",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"88",x"68",x"44",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"44",x"68",x"68",x"68",x"88",x"8c",x"ac",x"b0",x"d0",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"d0",x"88",x"40",x"40",x"20",x"20",x"20",x"44",x"68",x"68",x"68",x"68",x"88",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"8c",x"64",x"20",x"20",x"20",x"20",x"44",x"48",x"68",x"68",x"68",x"68",x"8c",x"8c",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f9",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"b0",x"ac",x"c8",x"c4",x"e0",x"c0",x"80",x"80",x"80",x"60",x"60",x"80",x"60",x"20",x"00",x"20",x"60",x"ad",x"d2"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"d2",x"ad",x"a9",x"84",x"80",x"60",x"60",x"64",x"69",x"6d",x"91",x"b1",x"d2",x"d2",x"f2",x"f2",x"f2",x"ed",x"e9",x"e9",x"e5",x"e5",x"e4",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"64",x"84",x"a4",x"c4",x"e4",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"40",x"20",x"20",x"20",x"40",x"40",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"84",x"ac",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f8",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fd",x"f8",x"fc",x"f8",x"f8",x"f8",x"f8",x"d0",x"cc",x"c4",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a8",x"ac",x"b0",x"d4",x"d4",x"f4",x"f9",x"fd",x"fd",x"fd",x"fd",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"b0",x"b0",x"8c",x"8c",x"88",x"64",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"40",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"44",x"64",x"68",x"68",x"88",x"8c",x"ac",x"b0",x"d0",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"d0",x"88",x"64",x"40",x"20",x"20",x"20",x"44",x"68",x"68",x"68",x"68",x"88",x"8c",x"8c",x"b0",x"d0",x"d0",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"ac",x"64",x"40",x"20",x"20",x"20",x"44",x"44",x"68",x"68",x"68",x"68",x"8c",x"8c",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f8",x"f4",x"f4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"b0",x"b0",x"ac",x"c4",x"e0",x"c0",x"80",x"80",x"80",x"60",x"60",x"80",x"60",x"20",x"00",x"20",x"60",x"ad",x"d2"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f7",x"d2",x"ad",x"a9",x"85",x"64",x"60",x"60",x"64",x"69",x"8d",x"8d",x"b1",x"b2",x"d2",x"d2",x"f2",x"f2",x"f2",x"ed",x"ed",x"e9",x"e5",x"e4",x"e4",x"e0",x"e4",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"60",x"64",x"84",x"84",x"a4",x"c4",x"c4",x"e4",x"e0",x"c0",x"a0",x"80",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"60",x"a8",x"f4",x"f4",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f8",x"d4",x"d4",x"d4",x"f4",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fd",x"fd",x"fe",x"fd",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"cc",x"c8",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"a0",x"80",x"80",x"a8",x"ac",x"d0",x"d0",x"d4",x"f8",x"f9",x"fd",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"8c",x"8c",x"88",x"64",x"40",x"40",x"60",x"60",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"64",x"68",x"68",x"88",x"8c",x"ac",x"b0",x"d0",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"ac",x"64",x"40",x"20",x"20",x"20",x"44",x"44",x"68",x"68",x"68",x"68",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"b0",x"68",x"44",x"20",x"20",x"20",x"40",x"44",x"68",x"68",x"68",x"68",x"8c",x"8c",x"b0",x"b0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f4",x"f4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"b0",x"ac",x"c8",x"e0",x"c0",x"80",x"80",x"80",x"60",x"60",x"80",x"60",x"20",x"00",x"20",x"60",x"ad",x"f2"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"d6",x"d2",x"ce",x"a9",x"84",x"60",x"60",x"40",x"40",x"64",x"69",x"91",x"b2",x"d6",x"d6",x"f6",x"f2",x"f2",x"ed",x"ed",x"ed",x"e9",x"e5",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"64",x"84",x"a4",x"a4",x"c4",x"c4",x"e4",x"c0",x"c0",x"a0",x"60",x"40",x"20",x"20",x"20",x"40",x"40",x"40",x"60",x"60",x"60",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"a8",x"d0",x"f4",x"d4",x"d4",x"d8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f8",x"d4",x"d4",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"cc",x"c4",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"a0",x"80",x"80",x"88",x"ac",x"d0",x"d0",x"d4",x"f4",x"f9",x"fd",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"8c",x"88",x"88",x"64",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"60",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"64",x"68",x"68",x"88",x"8c",x"ac",x"b0",x"d0",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"ac",x"88",x"44",x"20",x"20",x"20",x"40",x"44",x"64",x"68",x"68",x"68",x"88",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"b0",x"88",x"44",x"20",x"20",x"20",x"20",x"44",x"48",x"68",x"68",x"68",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f8",x"f4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"b0",x"90",x"c8",x"e0",x"c0",x"80",x"80",x"80",x"60",x"60",x"80",x"60",x"20",x"00",x"20",x"60",x"ad",x"f2"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"da",x"d2",x"ad",x"a9",x"84",x"80",x"60",x"60",x"64",x"89",x"89",x"8d",x"b2",x"b6",x"d6",x"f6",x"f6",x"f2",x"ee",x"ed",x"e9",x"e9",x"e9",x"e9",x"e5",x"e5",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"64",x"64",x"64",x"84",x"84",x"c4",x"c4",x"c4",x"c4",x"c0",x"a0",x"80",x"60",x"40",x"40",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"40",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"a4",x"cc",x"d4",x"d4",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f9",x"f9",x"f8",x"d4",x"d4",x"f8",x"fc",x"fc",x"fc",x"f8",x"fc",x"fd",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d0",x"b0",x"b0",x"b0",x"b0",x"b0",x"d0",x"d0",x"d0",x"d0",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"fd",x"fd",x"f9",x"f8",x"f8",x"f8",x"f8",x"f4",x"d0",x"cc",x"a4",x"a0",x"c0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"a0",x"80",x"a0",x"a0",x"88",x"ac",x"b0",x"d4",x"d0",x"f4",x"f9",x"fd",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"ac",x"88",x"64",x"60",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"64",x"68",x"68",x"88",x"8c",x"ac",x"b0",x"d0",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d0",x"b0",x"8c",x"64",x"40",x"20",x"20",x"40",x"44",x"44",x"68",x"68",x"68",x"68",x"8c",x"8c",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"8c",x"64",x"40",x"20",x"20",x"20",x"44",x"44",x"68",x"68",x"68",x"68",x"8c",x"ac",x"b0",x"b0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"fd",x"fd",x"fd",x"f9",x"f9",x"f8",x"f4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"b4",x"90",x"c8",x"e0",x"c0",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"20",x"00",x"20",x"60",x"cd",x"f6"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"db",x"d6",x"b2",x"ad",x"89",x"85",x"84",x"60",x"60",x"64",x"64",x"89",x"ad",x"b2",x"d6",x"f6",x"f6",x"f6",x"f2",x"f2",x"ed",x"e9",x"e9",x"e5",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"64",x"64",x"84",x"84",x"84",x"84",x"a4",x"a4",x"c4",x"e4",x"c4",x"c0",x"a0",x"80",x"60",x"40",x"20",x"00",x"00",x"00",x"20",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"84",x"cc",x"d0",x"d4",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f9",x"f8",x"d4",x"d8",x"f8",x"fc",x"fc",x"fc",x"f8",x"fc",x"fd",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"d4",x"d4",x"d0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"ac",x"ac",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"d0",x"d0",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d0",x"a8",x"a4",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"80",x"80",x"a0",x"a0",x"88",x"8c",x"b0",x"d0",x"d0",x"f4",x"f9",x"f9",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"ac",x"88",x"64",x"60",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"80",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"44",x"64",x"68",x"68",x"88",x"8c",x"ac",x"b0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d0",x"d0",x"ac",x"64",x"40",x"20",x"20",x"20",x"40",x"44",x"68",x"68",x"68",x"68",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"ac",x"68",x"40",x"20",x"20",x"20",x"20",x"44",x"68",x"68",x"68",x"68",x"8c",x"8c",x"b0",x"b0",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"fd",x"fd",x"fd",x"f9",x"f9",x"f9",x"f4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"d4",x"f4",x"f4",x"f4",x"d4",x"b4",x"b0",x"ac",x"c4",x"c0",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"20",x"00",x"20",x"60",x"ce",x"f6"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d2",x"ad",x"89",x"84",x"60",x"60",x"60",x"64",x"69",x"8d",x"91",x"b6",x"b6",x"d6",x"d6",x"f6",x"f6",x"f2",x"ee",x"ed",x"e9",x"e9",x"e9",x"e5",x"e4",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"84",x"84",x"a4",x"a4",x"c5",x"e5",x"e5",x"e5",x"c4",x"c0",x"c0",x"80",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"84",x"a8",x"d0",x"d4",x"d4",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f9",x"f8",x"f4",x"f8",x"fc",x"fc",x"fc",x"fc",x"fd",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"d4",x"b0",x"b0",x"b0",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"ac",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"fd",x"fd",x"fd",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"cc",x"a8",x"a4",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"a0",x"80",x"84",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f8",x"f9",x"fd",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"ac",x"88",x"64",x"60",x"60",x"60",x"60",x"60",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"44",x"64",x"68",x"68",x"8c",x"8c",x"b0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d0",x"d0",x"ac",x"68",x"40",x"40",x"20",x"20",x"20",x"44",x"68",x"68",x"68",x"68",x"88",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"88",x"44",x"20",x"20",x"20",x"20",x"44",x"68",x"68",x"68",x"68",x"8c",x"8c",x"b0",x"b0",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"fd",x"fd",x"fd",x"fd",x"f9",x"f9",x"f4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"d4",x"b4",x"b0",x"ac",x"c4",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"20",x"00",x"20",x"64",x"d2",x"f6"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"f7",x"d6",x"d2",x"cd",x"a9",x"84",x"60",x"60",x"60",x"64",x"89",x"8d",x"b2",x"b6",x"d6",x"da",x"fa",x"fa",x"f6",x"f2",x"ee",x"e9",x"e9",x"e5",x"e5",x"e4",x"e4",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"84",x"84",x"a4",x"a4",x"c4",x"e5",x"e5",x"e5",x"e4",x"c0",x"c0",x"a0",x"80",x"60",x"40",x"40",x"20",x"20",x"20",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"a8",x"d0",x"d4",x"d4",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f9",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"d4",x"b0",x"b0",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"6c",x"6c",x"6c",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"ac",x"b0",x"b0",x"b0",x"d0",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"fc",x"f8",x"f4",x"f4",x"f4",x"f4",x"f0",x"cc",x"a8",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"a0",x"80",x"84",x"8c",x"ac",x"ac",x"d0",x"d0",x"f4",x"f8",x"f9",x"fd",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"d0",x"b0",x"ac",x"88",x"64",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"44",x"64",x"68",x"88",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d0",x"d0",x"b0",x"88",x"44",x"40",x"20",x"20",x"20",x"44",x"68",x"68",x"68",x"68",x"68",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"b0",x"88",x"44",x"20",x"20",x"20",x"20",x"44",x"68",x"68",x"68",x"68",x"8c",x"8c",x"b0",x"b0",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"fd",x"fd",x"fd",x"fd",x"f9",x"f9",x"f4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"d4",x"d4",x"b0",x"ac",x"a4",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"20",x"00",x"20",x"64",x"d2",x"fb"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d7",x"b2",x"8e",x"89",x"80",x"60",x"60",x"64",x"64",x"69",x"8d",x"b2",x"d6",x"d6",x"f6",x"f6",x"f6",x"f6",x"f2",x"f2",x"ed",x"ed",x"e9",x"e5",x"e5",x"e5",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"84",x"84",x"84",x"a4",x"c4",x"e8",x"e9",x"e5",x"e4",x"e4",x"c0",x"a0",x"80",x"60",x"40",x"40",x"20",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"a4",x"ac",x"d4",x"d4",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f4",x"f4",x"f0",x"d0",x"ac",x"a4",x"a0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a4",x"88",x"8c",x"b0",x"d0",x"d0",x"f4",x"f4",x"f9",x"fd",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"d0",x"b0",x"ac",x"a8",x"64",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"44",x"64",x"68",x"88",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"88",x"64",x"40",x"20",x"20",x"20",x"44",x"68",x"68",x"68",x"68",x"68",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"b0",x"8c",x"44",x"20",x"20",x"20",x"20",x"44",x"68",x"68",x"68",x"68",x"8c",x"8c",x"b0",x"b0",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"fd",x"fd",x"fd",x"fd",x"f9",x"f9",x"f4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"d4",x"d4",x"b0",x"ac",x"a8",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"20",x"00",x"20",x"64",x"d2",x"fb"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f7",x"d6",x"b2",x"ad",x"89",x"69",x"64",x"60",x"64",x"64",x"89",x"8d",x"b2",x"b6",x"da",x"fa",x"fa",x"f6",x"f6",x"f2",x"ee",x"ed",x"e9",x"e5",x"e5",x"e4",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"64",x"64",x"64",x"64",x"84",x"84",x"a5",x"a4",x"c4",x"c4",x"c4",x"e4",x"e4",x"c4",x"c4",x"a0",x"80",x"60",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"84",x"ac",x"d4",x"d4",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"b0",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"68",x"68",x"68",x"68",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"ac",x"b0",x"b0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f5",x"f5",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"c8",x"a0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"80",x"84",x"88",x"8c",x"b0",x"b0",x"d0",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"d0",x"b0",x"ac",x"a8",x"84",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"44",x"64",x"68",x"8c",x"8c",x"b0",x"b0",x"d0",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"d0",x"8c",x"64",x"40",x"20",x"20",x"20",x"44",x"44",x"68",x"68",x"68",x"68",x"8c",x"8c",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"8c",x"64",x"40",x"20",x"20",x"20",x"44",x"68",x"68",x"68",x"68",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"fd",x"fd",x"fd",x"fd",x"f9",x"f9",x"f9",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d0",x"b0",x"ac",x"a4",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"20",x"20",x"40",x"84",x"d6",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"d2",x"ad",x"89",x"80",x"60",x"60",x"64",x"64",x"6d",x"92",x"92",x"b6",x"d6",x"fb",x"fb",x"fa",x"f6",x"f6",x"f2",x"ed",x"e9",x"e9",x"e9",x"e5",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"84",x"84",x"84",x"84",x"84",x"a4",x"c4",x"c5",x"e9",x"e5",x"e5",x"e4",x"c0",x"a0",x"80",x"60",x"40",x"40",x"20",x"20",x"40",x"40",x"40",x"60",x"60",x"40",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"60",x"88",x"d0",x"d4",x"d4",x"d4",x"f8",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"d4",x"d0",x"b0",x"8c",x"8c",x"8c",x"8c",x"6c",x"68",x"68",x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"68",x"6c",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"cc",x"c4",x"a0",x"a0",x"a0",x"a0",x"c0",x"a0",x"80",x"64",x"ac",x"ac",x"90",x"b0",x"d0",x"f0",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"d0",x"d0",x"d0",x"ac",x"84",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"44",x"64",x"68",x"8c",x"8c",x"b0",x"d0",x"d0",x"f4",x"f8",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"ac",x"88",x"40",x"20",x"20",x"20",x"40",x"44",x"68",x"68",x"68",x"68",x"88",x"8c",x"ac",x"b0",x"d0",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"ac",x"68",x"44",x"20",x"20",x"20",x"44",x"44",x"68",x"68",x"68",x"6c",x"8c",x"8c",x"b0",x"b0",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"f9",x"f9",x"f4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"d4",x"d4",x"b4",x"b4",x"b0",x"90",x"a8",x"a4",x"a0",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"20",x"20",x"60",x"84",x"f6",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"d2",x"d2",x"ad",x"a9",x"85",x"64",x"64",x"64",x"68",x"89",x"8d",x"b2",x"b6",x"da",x"da",x"fb",x"fa",x"f6",x"f6",x"f2",x"ed",x"e9",x"e9",x"e4",x"e4",x"e4",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"84",x"84",x"a4",x"a4",x"a4",x"a4",x"c4",x"c4",x"c4",x"c4",x"c4",x"c4",x"c0",x"a0",x"80",x"80",x"60",x"40",x"40",x"20",x"20",x"20",x"40",x"40",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"60",x"84",x"ac",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"d4",x"d0",x"b0",x"8c",x"8c",x"8c",x"6c",x"6c",x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"44",x"44",x"48",x"48",x"44",x"44",x"44",x"44",x"44",x"48",x"48",x"48",x"68",x"68",x"68",x"68",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d0",x"c8",x"a4",x"a0",x"a0",x"a0",x"c0",x"a0",x"80",x"84",x"88",x"8c",x"90",x"b0",x"d0",x"d0",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"d0",x"d0",x"d0",x"ac",x"84",x"60",x"60",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"44",x"64",x"68",x"8c",x"b0",x"b0",x"d0",x"d4",x"f4",x"f9",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"b0",x"88",x"64",x"20",x"20",x"20",x"40",x"44",x"68",x"68",x"68",x"68",x"68",x"8c",x"ac",x"b0",x"b0",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"b0",x"88",x"44",x"20",x"20",x"20",x"40",x"44",x"68",x"68",x"68",x"6c",x"8c",x"8c",x"b0",x"b0",x"d4",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"f9",x"f9",x"f4",x"f4",x"f4",x"f4",x"d4",x"f4",x"f4",x"f4",x"d4",x"b4",x"b0",x"b0",x"8c",x"88",x"a4",x"a0",x"80",x"80",x"80",x"80",x"60",x"40",x"40",x"20",x"20",x"60",x"a4",x"f6",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"da",x"d6",x"ad",x"a9",x"84",x"60",x"60",x"60",x"64",x"69",x"91",x"b6",x"b6",x"db",x"fb",x"fb",x"fa",x"fa",x"f6",x"f2",x"f2",x"ed",x"e9",x"e9",x"e9",x"e5",x"e5",x"e4",x"e0",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"64",x"64",x"84",x"84",x"84",x"84",x"a4",x"c5",x"e5",x"e5",x"e5",x"e5",x"e5",x"c4",x"a0",x"80",x"60",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"e0",x"e0",x"a0",x"a0",x"c0",x"c0",x"a0",x"80",x"60",x"84",x"ac",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"b0",x"8c",x"8c",x"8c",x"6c",x"68",x"48",x"48",x"48",x"48",x"48",x"44",x"64",x"64",x"64",x"64",x"64",x"44",x"64",x"64",x"44",x"44",x"64",x"64",x"44",x"44",x"64",x"68",x"68",x"68",x"68",x"68",x"8c",x"8c",x"8c",x"8c",x"ac",x"b0",x"b0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f0",x"cc",x"a4",x"a0",x"a0",x"c0",x"a0",x"a0",x"a0",x"84",x"88",x"8c",x"b0",x"b0",x"d0",x"d0",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"d0",x"d0",x"ac",x"84",x"60",x"60",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"a0",x"80",x"60",x"80",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"64",x"68",x"8c",x"b0",x"d0",x"d0",x"d4",x"f8",x"f9",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"b0",x"8c",x"64",x"20",x"20",x"40",x"40",x"40",x"44",x"68",x"68",x"68",x"68",x"8c",x"8c",x"b0",x"b0",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"b0",x"88",x"64",x"20",x"20",x"20",x"40",x"44",x"68",x"68",x"6c",x"6c",x"8c",x"8c",x"b0",x"b0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"fd",x"fd",x"fd",x"fd",x"f9",x"f9",x"f8",x"f4",x"f4",x"d4",x"d4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"90",x"8c",x"88",x"a4",x"a0",x"80",x"80",x"80",x"80",x"80",x"60",x"40",x"20",x"20",x"60",x"a5",x"f6",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"d2",x"b1",x"ad",x"89",x"89",x"84",x"64",x"64",x"64",x"89",x"8d",x"b2",x"b6",x"db",x"fb",x"fb",x"fb",x"f6",x"f6",x"f2",x"ed",x"ed",x"e9",x"e5",x"e5",x"e4",x"e4",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"84",x"84",x"84",x"a8",x"a9",x"a9",x"a9",x"c5",x"c5",x"e5",x"e5",x"c5",x"c4",x"a0",x"a0",x"80",x"60",x"60",x"40",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"64",x"84",x"84",x"a4",x"a4",x"a4",x"a4",x"a4",x"c4",x"c4",x"c4",x"c4",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"80",x"80",x"84",x"ac",x"d0",x"d4",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"b0",x"b0",x"8c",x"8c",x"88",x"68",x"68",x"68",x"48",x"48",x"48",x"44",x"44",x"64",x"64",x"64",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"44",x"44",x"64",x"64",x"64",x"64",x"64",x"68",x"8c",x"8c",x"8c",x"8c",x"8c",x"ac",x"b0",x"b0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f0",x"cc",x"a8",x"a4",x"a0",x"a0",x"a0",x"a0",x"a0",x"84",x"88",x"8c",x"8c",x"b0",x"b0",x"d0",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"d0",x"d0",x"ac",x"84",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"64",x"88",x"8c",x"b0",x"d0",x"d4",x"f4",x"f8",x"fd",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"ac",x"64",x"40",x"20",x"40",x"40",x"40",x"44",x"68",x"68",x"68",x"68",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"b0",x"8c",x"64",x"20",x"20",x"20",x"20",x"44",x"68",x"68",x"6c",x"6c",x"8c",x"8c",x"b0",x"b0",x"d4",x"d4",x"d4",x"f8",x"f8",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"fd",x"fd",x"fd",x"fd",x"f9",x"f9",x"f9",x"f4",x"f4",x"d4",x"d4",x"d4",x"f4",x"f4",x"d0",x"d0",x"b0",x"90",x"8c",x"88",x"a0",x"a0",x"80",x"80",x"60",x"80",x"80",x"60",x"20",x"20",x"20",x"60",x"a9",x"fb",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"ad",x"a8",x"80",x"60",x"60",x"60",x"64",x"89",x"8d",x"96",x"b6",x"da",x"fb",x"fb",x"fb",x"fb",x"f7",x"f2",x"ee",x"ed",x"e9",x"e9",x"e9",x"e5",x"e4",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"64",x"64",x"84",x"84",x"a8",x"a9",x"c9",x"e9",x"e9",x"e5",x"e5",x"e5",x"c5",x"a4",x"80",x"60",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"64",x"84",x"88",x"a8",x"a8",x"cc",x"cc",x"cc",x"cc",x"cc",x"ec",x"ec",x"ec",x"ec",x"ec",x"ec",x"e8",x"e8",x"c8",x"c8",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"e0",x"e0",x"c0",x"a0",x"e0",x"e0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"88",x"b0",x"d4",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"b0",x"90",x"8c",x"8c",x"68",x"68",x"68",x"68",x"48",x"44",x"44",x"44",x"44",x"64",x"60",x"60",x"60",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"60",x"60",x"44",x"44",x"64",x"64",x"64",x"64",x"68",x"68",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d0",x"d0",x"cc",x"c8",x"a0",x"a0",x"c0",x"a0",x"80",x"80",x"88",x"8c",x"8c",x"8c",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"d0",x"d0",x"ac",x"88",x"84",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"c0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"80",x"60",x"80",x"a0",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"68",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f8",x"fd",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"b0",x"68",x"40",x"40",x"40",x"40",x"40",x"44",x"48",x"68",x"68",x"68",x"8c",x"8c",x"ac",x"b0",x"d0",x"d0",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"d0",x"ac",x"64",x"20",x"20",x"20",x"20",x"44",x"68",x"6c",x"6c",x"6c",x"8c",x"8c",x"b0",x"b0",x"b0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"f9",x"f9",x"f4",x"f4",x"d4",x"d4",x"d4",x"f4",x"f0",x"d0",x"d0",x"b0",x"8c",x"8c",x"a8",x"a0",x"a0",x"80",x"60",x"60",x"80",x"80",x"60",x"20",x"20",x"40",x"84",x"c9",x"fb",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"f6",x"d2",x"d2",x"ad",x"89",x"88",x"84",x"64",x"64",x"89",x"89",x"ad",x"b2",x"d6",x"da",x"da",x"fb",x"fb",x"f6",x"f6",x"f2",x"ee",x"e9",x"e9",x"e5",x"e4",x"e4",x"e4",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"84",x"84",x"84",x"88",x"a8",x"a9",x"c9",x"c9",x"e5",x"e5",x"c5",x"c5",x"a4",x"a4",x"80",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"60",x"60",x"84",x"84",x"88",x"a8",x"a8",x"ac",x"cc",x"d0",x"d0",x"d0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"f0",x"ec",x"ec",x"e8",x"e8",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"84",x"ac",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"b0",x"90",x"8c",x"6c",x"6c",x"68",x"48",x"48",x"44",x"44",x"64",x"64",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"60",x"80",x"60",x"60",x"60",x"60",x"60",x"40",x"60",x"60",x"60",x"60",x"64",x"64",x"68",x"68",x"88",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"d0",x"cc",x"a4",x"a0",x"a0",x"a0",x"80",x"80",x"88",x"8c",x"8c",x"8c",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f4",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"d0",x"ac",x"a8",x"84",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"40",x"40",x"64",x"88",x"8c",x"b0",x"d0",x"d4",x"d4",x"f4",x"f9",x"fd",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"d0",x"88",x"40",x"40",x"40",x"40",x"40",x"44",x"44",x"68",x"68",x"68",x"88",x"8c",x"8c",x"b0",x"b0",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"68",x"40",x"20",x"20",x"20",x"44",x"48",x"68",x"6c",x"6c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"f9",x"f9",x"f9",x"f4",x"d4",x"d4",x"d4",x"d4",x"d0",x"d0",x"b0",x"ac",x"8c",x"88",x"a4",x"a0",x"a0",x"80",x"60",x"60",x"80",x"80",x"40",x"20",x"20",x"40",x"85",x"ce",x"fb",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"d6",x"ce",x"a9",x"a4",x"80",x"60",x"60",x"64",x"69",x"91",x"b6",x"db",x"fb",x"ff",x"ff",x"fb",x"fb",x"f6",x"f2",x"f2",x"ed",x"ed",x"e9",x"e5",x"e4",x"e4",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"84",x"84",x"84",x"a8",x"a9",x"c9",x"c9",x"e9",x"e9",x"e9",x"e5",x"c4",x"a0",x"80",x"60",x"40",x"20",x"20",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"64",x"88",x"ac",x"cc",x"d0",x"f4",x"f4",x"f4",x"f8",x"f9",x"f9",x"f9",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f0",x"ec",x"e8",x"e8",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"e0",x"e0",x"c0",x"c0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"84",x"ac",x"d0",x"d4",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"b0",x"b0",x"8c",x"6c",x"6c",x"68",x"48",x"48",x"44",x"44",x"64",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"44",x"64",x"68",x"68",x"88",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"cc",x"c4",x"a0",x"a0",x"80",x"a0",x"80",x"68",x"8c",x"8c",x"ac",x"b0",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"d0",x"ac",x"ac",x"84",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"60",x"80",x"a0",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"40",x"40",x"64",x"88",x"ac",x"d0",x"d0",x"d4",x"f4",x"f8",x"f9",x"fd",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"d0",x"88",x"64",x"40",x"40",x"20",x"20",x"40",x"44",x"68",x"68",x"68",x"68",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"b0",x"88",x"40",x"20",x"20",x"20",x"20",x"44",x"68",x"6c",x"6c",x"6c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f9",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"f9",x"f9",x"f9",x"f4",x"d4",x"d4",x"d4",x"d4",x"b0",x"b0",x"b0",x"8c",x"8c",x"a8",x"a4",x"a0",x"a0",x"80",x"60",x"60",x"80",x"80",x"40",x"20",x"20",x"40",x"a9",x"f2",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"d2",x"ad",x"a9",x"89",x"85",x"85",x"85",x"85",x"89",x"89",x"ae",x"b2",x"d6",x"db",x"db",x"fb",x"fb",x"fb",x"f6",x"f2",x"ee",x"ed",x"e9",x"e9",x"e5",x"e4",x"e4",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"84",x"84",x"a4",x"a5",x"a9",x"c9",x"c9",x"e9",x"e9",x"e5",x"c5",x"c4",x"a4",x"a4",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"00",x"00",x"20",x"20",x"00",x"00",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"64",x"88",x"88",x"ac",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f0",x"ec",x"e8",x"e8",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"a8",x"d0",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"8c",x"6c",x"6c",x"6c",x"68",x"48",x"44",x"44",x"64",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"44",x"64",x"68",x"68",x"88",x"8c",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"d0",x"c8",x"c0",x"80",x"80",x"a0",x"80",x"68",x"88",x"ac",x"ac",x"b0",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"d0",x"cc",x"a8",x"80",x"80",x"a0",x"a0",x"80",x"a0",x"a0",x"a0",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"40",x"40",x"64",x"ac",x"b0",x"d0",x"d4",x"d4",x"f4",x"f8",x"fd",x"fd",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"d0",x"ac",x"68",x"40",x"20",x"20",x"20",x"40",x"44",x"68",x"68",x"68",x"68",x"88",x"8c",x"ac",x"b0",x"b0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"8c",x"44",x"20",x"20",x"20",x"20",x"44",x"68",x"68",x"6c",x"6c",x"6c",x"8c",x"8c",x"8c",x"90",x"b0",x"b0",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f9",x"f9",x"f9",x"fd",x"fd",x"fd",x"f9",x"f9",x"f9",x"f5",x"d4",x"d4",x"d4",x"b4",x"b4",x"90",x"90",x"8c",x"8c",x"a8",x"a4",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"40",x"20",x"20",x"60",x"ad",x"f6",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fb",x"f7",x"f2",x"c9",x"a4",x"80",x"60",x"60",x"64",x"69",x"8d",x"b6",x"bb",x"db",x"fb",x"fb",x"fb",x"fb",x"f6",x"f6",x"f2",x"f2",x"ed",x"e9",x"e5",x"e5",x"e4",x"e4",x"e4",x"e4",x"c0",x"a0",x"a0",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"84",x"89",x"a9",x"c9",x"c9",x"e9",x"e9",x"e9",x"e5",x"e5",x"c4",x"a0",x"80",x"60",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"84",x"a8",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"f9",x"f8",x"f4",x"f0",x"ec",x"e4",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"e0",x"e0",x"c0",x"c0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"60",x"88",x"d0",x"d0",x"d4",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"b0",x"8c",x"8c",x"68",x"68",x"68",x"68",x"64",x"64",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"80",x"60",x"60",x"60",x"80",x"60",x"40",x"40",x"64",x"64",x"68",x"68",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"d0",x"c8",x"c4",x"80",x"80",x"a0",x"80",x"64",x"88",x"ac",x"ac",x"8c",x"b0",x"b0",x"d0",x"d0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"d0",x"d0",x"a8",x"84",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"a0",x"a0",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"60",x"80",x"80",x"60",x"60",x"40",x"40",x"64",x"88",x"ac",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"ac",x"88",x"44",x"20",x"20",x"20",x"20",x"44",x"68",x"68",x"68",x"68",x"88",x"8c",x"8c",x"b0",x"b0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"8c",x"64",x"40",x"20",x"20",x"20",x"44",x"44",x"68",x"68",x"68",x"6c",x"8c",x"8c",x"8c",x"8c",x"90",x"b0",x"b0",x"d0",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"d4",x"d4",x"d4",x"d0",x"b0",x"90",x"90",x"70",x"8c",x"88",x"a4",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"80",x"60",x"20",x"20",x"40",x"60",x"cd",x"fb",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"d2",x"ad",x"a9",x"a9",x"85",x"85",x"85",x"85",x"89",x"8d",x"91",x"b6",x"ba",x"db",x"fb",x"fb",x"fb",x"f7",x"f7",x"f2",x"ee",x"ed",x"e9",x"e9",x"e5",x"e5",x"e4",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"84",x"84",x"84",x"a4",x"a8",x"a9",x"c9",x"c9",x"c9",x"c9",x"c9",x"c5",x"c5",x"a4",x"a0",x"80",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"84",x"a8",x"cc",x"d0",x"f4",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f4",x"f0",x"f0",x"ec",x"e8",x"c4",x"c4",x"c0",x"c0",x"c0",x"e0",x"c0",x"c0",x"c0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"60",x"84",x"ac",x"d0",x"d4",x"d4",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"b0",x"b0",x"8c",x"8c",x"68",x"68",x"68",x"64",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"60",x"60",x"40",x"60",x"64",x"64",x"68",x"88",x"8c",x"8c",x"8c",x"ac",x"b0",x"b0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"d0",x"cc",x"a8",x"a0",x"80",x"80",x"80",x"84",x"88",x"8c",x"8c",x"8c",x"ac",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"d0",x"ac",x"a8",x"84",x"80",x"80",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"60",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"80",x"60",x"40",x"40",x"40",x"64",x"8c",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"b0",x"8c",x"64",x"20",x"20",x"20",x"20",x"40",x"44",x"68",x"68",x"68",x"8c",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"ac",x"68",x"44",x"20",x"20",x"20",x"20",x"44",x"44",x"68",x"68",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"90",x"b0",x"b0",x"b0",x"b0",x"b0",x"d0",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d9",x"d9",x"f9",x"d5",x"d5",x"d4",x"d4",x"d0",x"b0",x"b0",x"90",x"90",x"70",x"6c",x"8c",x"a8",x"c4",x"e0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"60",x"40",x"20",x"20",x"40",x"80",x"d2",x"fb",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"d2",x"ad",x"89",x"64",x"60",x"40",x"60",x"89",x"8e",x"b2",x"b6",x"db",x"df",x"ff",x"ff",x"fb",x"fa",x"f6",x"f2",x"ed",x"ed",x"ed",x"e9",x"e4",x"e4",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"84",x"84",x"84",x"84",x"a8",x"a9",x"c9",x"cd",x"c9",x"e9",x"e9",x"e9",x"c5",x"c4",x"a4",x"80",x"40",x"40",x"20",x"20",x"40",x"40",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"a4",x"ac",x"d0",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fc",x"f8",x"f8",x"fc",x"f8",x"f8",x"f8",x"f4",x"f4",x"f0",x"ec",x"cc",x"c4",x"c0",x"e0",x"e0",x"c0",x"a0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"84",x"a8",x"b0",x"d0",x"d4",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f8",x"f9",x"f9",x"f9",x"d4",x"b0",x"b0",x"8c",x"8c",x"88",x"68",x"68",x"64",x"64",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"64",x"64",x"68",x"88",x"8c",x"8c",x"8c",x"ac",x"b0",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"d0",x"cc",x"a8",x"a0",x"80",x"80",x"60",x"84",x"88",x"8c",x"8c",x"8c",x"ac",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"cc",x"a8",x"a4",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"60",x"60",x"a0",x"a0",x"80",x"60",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"60",x"60",x"60",x"40",x"64",x"88",x"ac",x"d0",x"f4",x"f4",x"f4",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"d0",x"ac",x"64",x"40",x"20",x"20",x"20",x"20",x"44",x"68",x"68",x"68",x"8c",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"b0",x"88",x"44",x"20",x"20",x"20",x"20",x"20",x"44",x"44",x"68",x"6c",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"d0",x"d0",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d0",x"b0",x"b0",x"b0",x"90",x"90",x"70",x"6c",x"6c",x"88",x"a4",x"c0",x"e0",x"c0",x"80",x"80",x"80",x"80",x"80",x"60",x"40",x"20",x"20",x"40",x"84",x"d2",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"d2",x"ad",x"a9",x"89",x"85",x"85",x"85",x"89",x"89",x"8d",x"92",x"b6",x"bb",x"db",x"db",x"fb",x"fb",x"f6",x"f6",x"f2",x"f2",x"ed",x"ed",x"e9",x"e8",x"e4",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"80",x"84",x"84",x"84",x"a5",x"a9",x"a9",x"a9",x"c9",x"c9",x"c9",x"c9",x"c9",x"c5",x"c4",x"a4",x"a4",x"80",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"84",x"a4",x"ac",x"d0",x"f4",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"ec",x"e8",x"c4",x"c4",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"88",x"ac",x"d0",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f8",x"f9",x"f9",x"f9",x"d4",x"b0",x"8c",x"8c",x"8c",x"88",x"88",x"64",x"64",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"64",x"64",x"68",x"88",x"8c",x"8c",x"ac",x"ac",x"b0",x"b0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"d0",x"d0",x"cc",x"a4",x"80",x"80",x"80",x"60",x"64",x"8c",x"8c",x"8c",x"8c",x"ac",x"b0",x"d0",x"d0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"d0",x"cc",x"a8",x"84",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"60",x"60",x"60",x"64",x"68",x"8c",x"d0",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"68",x"40",x"20",x"20",x"20",x"20",x"40",x"44",x"68",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"b0",x"8c",x"64",x"20",x"20",x"20",x"20",x"20",x"20",x"44",x"48",x"68",x"68",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"90",x"90",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"88",x"a4",x"c4",x"c0",x"e0",x"c0",x"80",x"80",x"80",x"80",x"80",x"60",x"40",x"20",x"20",x"60",x"a5",x"d6",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fa",x"d2",x"ad",x"89",x"80",x"60",x"60",x"60",x"64",x"89",x"b2",x"b6",x"da",x"df",x"df",x"df",x"ff",x"fb",x"f6",x"f2",x"ee",x"ed",x"e9",x"e9",x"e8",x"e4",x"e4",x"e0",x"e0",x"e0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"64",x"84",x"84",x"84",x"84",x"a4",x"a9",x"a9",x"c9",x"cd",x"cd",x"e9",x"e9",x"c9",x"c5",x"c4",x"a0",x"80",x"60",x"40",x"40",x"20",x"20",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"a4",x"a8",x"d0",x"f4",x"f9",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"f8",x"f4",x"ec",x"cc",x"a8",x"c4",x"c0",x"c0",x"a0",x"c0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"84",x"ac",x"d0",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f9",x"f9",x"d4",x"b4",x"90",x"8c",x"6c",x"88",x"88",x"84",x"64",x"60",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"60",x"60",x"60",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"64",x"68",x"88",x"8c",x"8c",x"ac",x"ac",x"ac",x"b0",x"d0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"f0",x"cc",x"a4",x"80",x"80",x"80",x"40",x"64",x"88",x"8c",x"8c",x"8c",x"ac",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"d0",x"d0",x"cc",x"a4",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"a0",x"80",x"60",x"60",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"40",x"60",x"80",x"60",x"60",x"60",x"60",x"60",x"64",x"68",x"8c",x"b0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"b0",x"88",x"44",x"40",x"20",x"20",x"20",x"40",x"44",x"68",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"8c",x"64",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"44",x"48",x"68",x"68",x"6c",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"90",x"90",x"90",x"90",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"6c",x"8c",x"a8",x"a4",x"c4",x"c0",x"e0",x"e0",x"a0",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"20",x"20",x"80",x"c9",x"f6",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"b2",x"ad",x"a9",x"89",x"84",x"64",x"64",x"69",x"89",x"8d",x"b2",x"d6",x"d6",x"db",x"fb",x"fb",x"fb",x"f6",x"f6",x"f6",x"f2",x"ed",x"e9",x"e9",x"e5",x"e4",x"e4",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"84",x"84",x"88",x"88",x"a8",x"a9",x"c9",x"c9",x"e9",x"e9",x"e9",x"e9",x"c4",x"a4",x"84",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"84",x"a8",x"cc",x"f0",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f0",x"cc",x"c8",x"c4",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"84",x"ac",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f9",x"f9",x"d4",x"b0",x"90",x"8c",x"6c",x"68",x"88",x"84",x"64",x"60",x"60",x"60",x"80",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"80",x"60",x"60",x"60",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"64",x"64",x"68",x"88",x"8c",x"8c",x"ac",x"ac",x"b0",x"d0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"d0",x"d0",x"cc",x"c8",x"a0",x"60",x"60",x"60",x"64",x"68",x"88",x"8c",x"ac",x"ac",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f4",x"d4",x"d4",x"d4",x"d4",x"f0",x"cc",x"a4",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"60",x"60",x"60",x"80",x"60",x"60",x"60",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"64",x"88",x"ac",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"b0",x"8c",x"64",x"40",x"20",x"20",x"20",x"20",x"44",x"68",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f8",x"f4",x"d4",x"f4",x"f4",x"f4",x"d4",x"d0",x"ac",x"64",x"20",x"20",x"20",x"20",x"00",x"20",x"20",x"20",x"24",x"44",x"68",x"68",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"b0",x"90",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"6c",x"6c",x"88",x"a4",x"c0",x"e0",x"e0",x"e0",x"e0",x"a0",x"60",x"80",x"80",x"80",x"60",x"40",x"40",x"20",x"20",x"80",x"c9",x"fb",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"b2",x"8e",x"89",x"64",x"60",x"60",x"60",x"64",x"69",x"91",x"b6",x"da",x"ff",x"ff",x"ff",x"fb",x"fb",x"f6",x"f2",x"ed",x"ed",x"e9",x"e9",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"60",x"64",x"84",x"84",x"84",x"a8",x"a9",x"a9",x"a8",x"a9",x"c9",x"c9",x"e9",x"e9",x"e5",x"c4",x"a0",x"80",x"60",x"40",x"40",x"20",x"20",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a4",x"a8",x"d0",x"f4",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"cc",x"c8",x"c4",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"84",x"ac",x"d0",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"b0",x"90",x"8c",x"68",x"68",x"88",x"84",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"64",x"64",x"88",x"8c",x"8c",x"ac",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"d0",x"b0",x"ac",x"c8",x"a4",x"60",x"40",x"60",x"64",x"44",x"68",x"8c",x"ac",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"d4",x"f4",x"f4",x"cc",x"a8",x"84",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"60",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"88",x"ac",x"b0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"b0",x"8c",x"68",x"40",x"20",x"20",x"20",x"20",x"40",x"68",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f8",x"f4",x"d4",x"f4",x"f4",x"f4",x"d4",x"d4",x"ac",x"64",x"20",x"20",x"20",x"20",x"00",x"20",x"20",x"20",x"20",x"24",x"44",x"48",x"68",x"6c",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"ac",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"6c",x"6c",x"88",x"a8",x"c4",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"60",x"80",x"80",x"80",x"60",x"40",x"40",x"20",x"40",x"a4",x"ee",x"fb",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"d2",x"ad",x"89",x"85",x"64",x"64",x"65",x"69",x"89",x"8d",x"8d",x"b2",x"d6",x"da",x"fa",x"fa",x"fa",x"f6",x"f6",x"f2",x"ed",x"ed",x"e9",x"e9",x"e5",x"e4",x"e4",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"84",x"84",x"84",x"a9",x"a9",x"c9",x"c9",x"e9",x"e9",x"e9",x"c9",x"c8",x"a4",x"84",x"80",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"c8",x"cc",x"f4",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"f9",x"f8",x"f8",x"f8",x"f8",x"d4",x"d0",x"cc",x"c4",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"a8",x"d0",x"d0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f5",x"f5",x"f4",x"d4",x"b4",x"90",x"8c",x"8c",x"88",x"68",x"64",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"60",x"60",x"60",x"80",x"60",x"60",x"60",x"64",x"64",x"88",x"8c",x"ac",x"ac",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"d0",x"d0",x"cc",x"cc",x"a4",x"60",x"60",x"60",x"60",x"64",x"68",x"8c",x"8c",x"8c",x"ac",x"ac",x"b0",x"d0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"cc",x"a8",x"84",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"60",x"60",x"84",x"ac",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"d0",x"ac",x"88",x"40",x"20",x"20",x"20",x"20",x"40",x"68",x"68",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"b0",x"88",x"40",x"20",x"20",x"20",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"24",x"44",x"48",x"68",x"68",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"ac",x"8c",x"90",x"70",x"6c",x"6c",x"8c",x"8c",x"8c",x"8c",x"6c",x"6c",x"68",x"88",x"a8",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"80",x"80",x"60",x"60",x"80",x"80",x"40",x"20",x"40",x"80",x"cd",x"f6",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"fa",x"d2",x"cd",x"a9",x"84",x"60",x"60",x"60",x"64",x"89",x"92",x"b6",x"d6",x"db",x"fb",x"fb",x"fb",x"fa",x"f6",x"f2",x"ed",x"ed",x"e9",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"64",x"84",x"84",x"84",x"84",x"84",x"84",x"a4",x"a8",x"a9",x"a9",x"c9",x"c9",x"e9",x"e9",x"e9",x"e9",x"e9",x"c5",x"a4",x"80",x"60",x"40",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"c0",x"c0",x"a0",x"c4",x"ec",x"f4",x"f8",x"fc",x"fc",x"fc",x"fd",x"fc",x"fc",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"f9",x"f8",x"f8",x"fc",x"d8",x"d8",x"d0",x"cc",x"c4",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"60",x"84",x"cc",x"d0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f9",x"f5",x"d4",x"d4",x"b0",x"90",x"8c",x"88",x"88",x"84",x"64",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"60",x"60",x"60",x"60",x"64",x"88",x"88",x"8c",x"ac",x"b0",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"d0",x"d0",x"cc",x"ac",x"a8",x"80",x"60",x"60",x"60",x"64",x"68",x"68",x"8c",x"8c",x"8c",x"8c",x"ac",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"d0",x"ac",x"88",x"64",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"80",x"80",x"60",x"64",x"a8",x"d0",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fd",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"d0",x"d0",x"ac",x"64",x"20",x"20",x"20",x"20",x"20",x"44",x"68",x"6c",x"8c",x"8c",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"8c",x"64",x"40",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"24",x"44",x"48",x"48",x"68",x"6c",x"6c",x"6c",x"6c",x"8c",x"8c",x"8c",x"90",x"70",x"6c",x"68",x"68",x"88",x"8c",x"6c",x"6c",x"69",x"69",x"a8",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"60",x"60",x"60",x"80",x"40",x"20",x"60",x"a0",x"f2",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"d2",x"a9",x"85",x"84",x"84",x"64",x"64",x"69",x"8d",x"b1",x"b6",x"d6",x"da",x"fb",x"fa",x"f6",x"f6",x"f2",x"f2",x"ee",x"ed",x"e9",x"e9",x"e5",x"e4",x"e4",x"e4",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"84",x"84",x"84",x"84",x"88",x"89",x"8d",x"ad",x"cd",x"ed",x"e9",x"e9",x"e9",x"c5",x"c4",x"a4",x"84",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c8",x"ec",x"f0",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"f9",x"f8",x"f8",x"f4",x"f4",x"d0",x"cc",x"c8",x"c0",x"c0",x"c0",x"c0",x"e0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"60",x"84",x"a8",x"d0",x"d0",x"d4",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f5",x"f4",x"d4",x"b4",x"b0",x"b0",x"8c",x"8c",x"88",x"84",x"80",x"60",x"60",x"80",x"80",x"60",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"64",x"84",x"88",x"8c",x"ac",x"b0",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"d0",x"d0",x"cc",x"ac",x"a8",x"80",x"60",x"60",x"60",x"64",x"64",x"68",x"8c",x"8c",x"8c",x"8c",x"ac",x"b0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"cc",x"ac",x"88",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"84",x"88",x"cc",x"d0",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"d0",x"ac",x"64",x"40",x"20",x"20",x"20",x"20",x"44",x"68",x"6c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"d0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"8c",x"64",x"40",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"24",x"24",x"44",x"48",x"48",x"48",x"48",x"68",x"88",x"88",x"6c",x"68",x"48",x"48",x"68",x"88",x"88",x"68",x"48",x"48",x"69",x"c4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"60",x"60",x"60",x"60",x"40",x"40",x"60",x"a0",x"f2",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d2",x"ad",x"85",x"80",x"60",x"60",x"64",x"89",x"8d",x"b2",x"b6",x"da",x"fb",x"fb",x"fb",x"fa",x"f6",x"f2",x"ed",x"ed",x"e9",x"e5",x"e5",x"e4",x"e4",x"e4",x"c0",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"84",x"a4",x"a4",x"a4",x"a4",x"a9",x"a9",x"ad",x"ad",x"cd",x"cd",x"e9",x"e9",x"e5",x"c4",x"a0",x"80",x"80",x"40",x"20",x"20",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"a0",x"80",x"80",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"a0",x"c4",x"f0",x"f5",x"f5",x"f8",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"fd",x"f9",x"f8",x"f4",x"f4",x"f8",x"f4",x"d4",x"cc",x"c4",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"84",x"a8",x"ac",x"d0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f5",x"f4",x"d4",x"b0",x"b0",x"90",x"8c",x"88",x"88",x"84",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"80",x"60",x"60",x"64",x"84",x"88",x"8c",x"ac",x"b0",x"b0",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"d0",x"d0",x"d0",x"ac",x"a8",x"80",x"60",x"60",x"60",x"60",x"64",x"68",x"8c",x"8c",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"d0",x"ac",x"84",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"80",x"60",x"80",x"a8",x"d0",x"d0",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"d0",x"ac",x"64",x"40",x"40",x"20",x"20",x"20",x"44",x"68",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"ac",x"68",x"40",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"24",x"24",x"24",x"24",x"44",x"64",x"64",x"64",x"44",x"44",x"44",x"64",x"84",x"84",x"44",x"48",x"48",x"68",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"60",x"40",x"40",x"60",x"80",x"a5",x"f2",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"ce",x"a5",x"84",x"60",x"64",x"64",x"69",x"8d",x"b2",x"d6",x"da",x"fb",x"fb",x"f6",x"f6",x"f2",x"f2",x"ed",x"ed",x"e9",x"e9",x"e5",x"e4",x"e4",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"84",x"84",x"88",x"89",x"ad",x"cd",x"ed",x"ed",x"e9",x"e9",x"e5",x"c4",x"a4",x"60",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c8",x"cc",x"f5",x"f9",x"f9",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fd",x"f9",x"f8",x"f8",x"f8",x"f8",x"f4",x"f0",x"ec",x"c8",x"c4",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"84",x"ac",x"d0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f5",x"f4",x"d4",x"b0",x"b0",x"90",x"8c",x"88",x"84",x"64",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"64",x"88",x"8c",x"8c",x"ac",x"b0",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"d0",x"d0",x"ac",x"a8",x"84",x"60",x"60",x"60",x"60",x"64",x"68",x"68",x"8c",x"8c",x"8c",x"8c",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d0",x"a8",x"84",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"80",x"84",x"a8",x"d0",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"b0",x"88",x"64",x"40",x"20",x"20",x"20",x"40",x"44",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"d4",x"d4",x"d4",x"f8",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"b0",x"88",x"44",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"24",x"24",x"48",x"88",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"80",x"40",x"20",x"60",x"80",x"a4",x"c9",x"f6",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b2",x"a9",x"a5",x"80",x"60",x"60",x"65",x"8d",x"b2",x"d6",x"fa",x"fb",x"fb",x"f6",x"f2",x"f2",x"ed",x"e9",x"e9",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"84",x"84",x"84",x"84",x"84",x"88",x"a9",x"a9",x"a9",x"a9",x"cd",x"ed",x"ed",x"e9",x"e5",x"c5",x"c0",x"a0",x"60",x"40",x"20",x"20",x"20",x"40",x"40",x"60",x"80",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"40",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"c0",x"c4",x"ec",x"f4",x"f8",x"fd",x"fc",x"fc",x"fc",x"fd",x"fd",x"fe",x"fe",x"fe",x"ff",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fd",x"f9",x"f9",x"f8",x"f8",x"f8",x"f4",x"f0",x"cc",x"c8",x"c4",x"a0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"64",x"a8",x"d0",x"d0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f5",x"f4",x"d0",x"b0",x"90",x"8c",x"8c",x"88",x"84",x"64",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"a0",x"c0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"64",x"88",x"8c",x"8c",x"ac",x"b0",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"d0",x"b0",x"ac",x"a8",x"84",x"60",x"60",x"60",x"60",x"64",x"64",x"68",x"8c",x"8c",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d0",x"ac",x"a8",x"a4",x"80",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"84",x"a8",x"cc",x"f0",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"b0",x"8c",x"64",x"40",x"20",x"40",x"20",x"20",x"44",x"68",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"d0",x"d4",x"d4",x"f8",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"f9",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"b0",x"8c",x"44",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"40",x"40",x"40",x"40",x"40",x"60",x"80",x"60",x"40",x"24",x"24",x"64",x"a4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"40",x"20",x"60",x"a0",x"c5",x"ce",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"f6",x"ce",x"89",x"64",x"40",x"44",x"69",x"8d",x"b1",x"d2",x"d6",x"f6",x"f6",x"f6",x"f2",x"ee",x"e9",x"e9",x"e5",x"e5",x"e5",x"e4",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"84",x"84",x"84",x"88",x"89",x"ad",x"ad",x"cd",x"ed",x"ed",x"e9",x"e5",x"c5",x"a4",x"80",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e4",x"ec",x"f4",x"f8",x"f8",x"fc",x"fc",x"fc",x"fd",x"fd",x"fe",x"ff",x"ff",x"ff",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fd",x"f9",x"f8",x"f4",x"f4",x"f4",x"d4",x"cc",x"c8",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"60",x"60",x"88",x"ac",x"b0",x"b0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f5",x"d4",x"b0",x"b0",x"8c",x"8c",x"8c",x"88",x"64",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"c0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"c0",x"c0",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"64",x"88",x"a8",x"8c",x"ac",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"d0",x"b0",x"b0",x"ac",x"84",x"60",x"60",x"60",x"40",x"40",x"44",x"68",x"68",x"8c",x"8c",x"8c",x"ac",x"b0",x"b0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d0",x"cc",x"a8",x"84",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"84",x"88",x"ac",x"d0",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f9",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"ac",x"88",x"40",x"40",x"40",x"20",x"20",x"40",x"68",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"d4",x"d4",x"f8",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"f9",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"ac",x"64",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"80",x"80",x"60",x"20",x"04",x"24",x"84",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"80",x"60",x"60",x"80",x"80",x"80",x"40",x"20",x"80",x"c0",x"c9",x"f6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"ad",x"85",x"60",x"60",x"44",x"48",x"91",x"d6",x"d6",x"f6",x"f6",x"f6",x"f2",x"ed",x"e9",x"e5",x"e5",x"e4",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"84",x"84",x"84",x"89",x"a9",x"a9",x"a9",x"ad",x"cd",x"cd",x"cd",x"c9",x"c9",x"c5",x"c0",x"a0",x"80",x"40",x"20",x"20",x"20",x"20",x"40",x"60",x"80",x"80",x"80",x"60",x"60",x"40",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e4",x"ec",x"f4",x"f8",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fe",x"ff",x"ff",x"ff",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"f5",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fd",x"f8",x"f8",x"f4",x"f8",x"d4",x"d0",x"cc",x"c8",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"60",x"60",x"88",x"ac",x"b0",x"d0",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"b0",x"b0",x"8c",x"8c",x"8c",x"88",x"64",x"80",x"80",x"60",x"60",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"a0",x"c0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"c0",x"a0",x"80",x"a0",x"a0",x"80",x"60",x"60",x"80",x"60",x"60",x"60",x"60",x"84",x"88",x"8c",x"ac",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"b0",x"ac",x"84",x"60",x"60",x"60",x"40",x"40",x"44",x"64",x"68",x"8c",x"8c",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"cc",x"a8",x"a8",x"84",x"84",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"84",x"84",x"a8",x"cc",x"d0",x"f4",x"f8",x"f8",x"f8",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"d0",x"ac",x"88",x"60",x"40",x"40",x"20",x"20",x"40",x"68",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"d4",x"d4",x"f8",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"f9",x"f9",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"b0",x"64",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"40",x"40",x"20",x"40",x"60",x"80",x"80",x"40",x"04",x"05",x"45",x"c4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"60",x"80",x"80",x"60",x"40",x"40",x"80",x"c0",x"ed",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"d6",x"a9",x"84",x"60",x"60",x"64",x"89",x"b1",x"d2",x"d6",x"f6",x"f2",x"f1",x"ed",x"e9",x"e9",x"e5",x"e5",x"e5",x"e4",x"e4",x"c0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"80",x"84",x"84",x"80",x"80",x"84",x"89",x"a9",x"ad",x"cd",x"cd",x"ed",x"ed",x"e9",x"e9",x"e9",x"c5",x"a4",x"84",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"48",x"48",x"48",x"48",x"48",x"44",x"44",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"60",x"60",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e8",x"f0",x"f8",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fe",x"ff",x"ff",x"ff",x"fe",x"fd",x"fd",x"fc",x"fc",x"fc",x"fd",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d0",x"d0",x"d0",x"d0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"d0",x"d4",x"d4",x"d4",x"d4",x"f5",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"fd",x"fd",x"fe",x"fe",x"fe",x"fd",x"fd",x"f8",x"f8",x"f4",x"d4",x"d0",x"d0",x"cc",x"c8",x"c0",x"c0",x"a0",x"c0",x"c0",x"a0",x"80",x"60",x"80",x"84",x"8c",x"b0",x"d0",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d0",x"b0",x"b0",x"8c",x"8c",x"8c",x"88",x"84",x"60",x"60",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"e0",x"c0",x"a0",x"c0",x"e0",x"c0",x"a0",x"c0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"c0",x"a0",x"a0",x"e0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"64",x"88",x"ac",x"ac",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"b0",x"ac",x"84",x"60",x"60",x"60",x"40",x"40",x"40",x"44",x"68",x"68",x"8c",x"8c",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f0",x"cc",x"cc",x"a8",x"84",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"84",x"ac",x"d0",x"f0",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f9",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"8c",x"64",x"40",x"40",x"20",x"20",x"40",x"64",x"68",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"b0",x"d4",x"d4",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"f9",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"d4",x"b0",x"68",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"40",x"40",x"20",x"20",x"60",x"80",x"80",x"80",x"20",x"04",x"25",x"65",x"c4",x"e0",x"e4",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"80",x"80",x"60",x"40",x"40",x"60",x"80",x"c4",x"f2",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d2",x"a9",x"80",x"60",x"60",x"60",x"89",x"d1",x"f2",x"f6",x"f2",x"ed",x"ed",x"e9",x"e5",x"e4",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"60",x"60",x"80",x"60",x"60",x"60",x"60",x"60",x"80",x"84",x"84",x"84",x"84",x"a4",x"a4",x"a4",x"a9",x"c9",x"cd",x"cd",x"ed",x"ed",x"ed",x"e9",x"c9",x"c5",x"a4",x"a0",x"80",x"60",x"40",x"20",x"20",x"40",x"60",x"60",x"80",x"80",x"80",x"60",x"40",x"40",x"20",x"20",x"20",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"20",x"24",x"24",x"48",x"6c",x"90",x"90",x"90",x"b0",x"b0",x"90",x"8c",x"88",x"84",x"84",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"e0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e4",x"e8",x"f0",x"f4",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fe",x"ff",x"ff",x"ff",x"fe",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"d4",x"d4",x"d0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"90",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"d0",x"d4",x"d4",x"d4",x"d5",x"f5",x"f5",x"f5",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"fe",x"fe",x"fe",x"fd",x"fd",x"f8",x"f4",x"f4",x"f0",x"d0",x"d0",x"cc",x"c4",x"c0",x"a0",x"a0",x"c0",x"a0",x"80",x"80",x"60",x"84",x"88",x"ac",x"d0",x"d0",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d0",x"b0",x"b0",x"8c",x"8c",x"8c",x"84",x"80",x"60",x"60",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"a0",x"c0",x"e0",x"c0",x"a0",x"c0",x"e0",x"c0",x"c0",x"c0",x"e0",x"c0",x"c0",x"c0",x"c0",x"e0",x"c0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"64",x"88",x"ac",x"ac",x"b0",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"b0",x"ac",x"84",x"60",x"60",x"60",x"40",x"40",x"40",x"44",x"64",x"68",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f0",x"d0",x"ac",x"a8",x"a4",x"84",x"84",x"84",x"84",x"84",x"84",x"88",x"a8",x"cc",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f8",x"f8",x"f4",x"d4",x"d4",x"d4",x"b0",x"8c",x"64",x"40",x"40",x"40",x"20",x"40",x"44",x"68",x"8c",x"8c",x"8c",x"8c",x"90",x"b0",x"b0",x"b0",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"f9",x"f9",x"f4",x"d4",x"d4",x"d4",x"d4",x"d4",x"b0",x"68",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"40",x"40",x"20",x"20",x"60",x"a0",x"80",x"60",x"04",x"04",x"45",x"a5",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"60",x"80",x"80",x"60",x"40",x"60",x"80",x"a0",x"c9",x"f6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"f6",x"cd",x"84",x"60",x"40",x"44",x"89",x"cd",x"ed",x"ed",x"ed",x"ed",x"e9",x"e5",x"e5",x"e4",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"84",x"84",x"a9",x"a9",x"a9",x"cd",x"cd",x"ed",x"e9",x"e9",x"e9",x"e9",x"c5",x"a4",x"60",x"40",x"20",x"20",x"20",x"40",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"68",x"ac",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"d4",x"d0",x"cc",x"a8",x"a4",x"80",x"80",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e4",x"ec",x"f4",x"f8",x"fc",x"fc",x"fc",x"fd",x"fd",x"fe",x"ff",x"ff",x"ff",x"fe",x"fd",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"d4",x"d0",x"b0",x"b0",x"b0",x"b0",x"ac",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"b0",x"d0",x"d4",x"d4",x"f4",x"f5",x"f9",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fe",x"fd",x"fd",x"f9",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"c8",x"c4",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"60",x"80",x"a4",x"ac",x"b0",x"d0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d0",x"b0",x"b0",x"ac",x"ac",x"88",x"88",x"64",x"80",x"80",x"80",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"c0",x"e0",x"c0",x"a0",x"c0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"c0",x"a0",x"a0",x"e0",x"c0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"60",x"60",x"80",x"80",x"40",x"40",x"84",x"a8",x"ac",x"b0",x"b0",x"d0",x"d0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"b0",x"ac",x"84",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"44",x"68",x"88",x"8c",x"8c",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f0",x"f0",x"f0",x"d0",x"f0",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f8",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"fd",x"f9",x"f9",x"f8",x"f8",x"f8",x"d4",x"d4",x"d4",x"b0",x"ac",x"64",x"40",x"40",x"40",x"20",x"40",x"40",x"64",x"88",x"8c",x"8c",x"8c",x"90",x"b0",x"b0",x"b0",x"d4",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"f9",x"f9",x"f4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d0",x"88",x"44",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"40",x"40",x"20",x"40",x"80",x"a0",x"60",x"20",x"04",x"04",x"84",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"40",x"60",x"a0",x"a4",x"cd",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fa",x"d2",x"a9",x"84",x"60",x"60",x"64",x"89",x"ad",x"ed",x"ed",x"e9",x"e9",x"e5",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"84",x"84",x"84",x"89",x"a9",x"a9",x"a9",x"c9",x"c9",x"cd",x"ed",x"e9",x"c9",x"c5",x"c5",x"a4",x"80",x"60",x"40",x"40",x"20",x"20",x"20",x"40",x"60",x"80",x"80",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"44",x"68",x"b0",x"f4",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"f9",x"f4",x"d0",x"cc",x"a8",x"84",x"a4",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c4",x"e8",x"f4",x"f9",x"fd",x"fc",x"fc",x"fc",x"fd",x"fe",x"ff",x"ff",x"ff",x"fe",x"fd",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"d4",x"d0",x"b0",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"6c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"b0",x"d0",x"d4",x"d4",x"f5",x"f9",x"f9",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"f8",x"f4",x"f4",x"d4",x"d4",x"d0",x"cc",x"c4",x"c4",x"a0",x"a0",x"a0",x"a0",x"80",x"60",x"80",x"84",x"ac",x"b0",x"d0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d0",x"b0",x"b0",x"ac",x"ac",x"88",x"88",x"64",x"80",x"80",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"c0",x"a0",x"c0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"c0",x"a0",x"c0",x"e0",x"c0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"60",x"80",x"60",x"40",x"40",x"84",x"88",x"ac",x"b0",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"b0",x"ac",x"84",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"44",x"64",x"68",x"88",x"8c",x"8c",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"fd",x"fd",x"f9",x"f9",x"f8",x"d4",x"d4",x"d4",x"d4",x"b0",x"8c",x"64",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"68",x"8c",x"8c",x"8c",x"90",x"b0",x"b0",x"b0",x"d4",x"d4",x"d4",x"f8",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"f9",x"f9",x"f8",x"d4",x"f8",x"d4",x"d4",x"d4",x"d4",x"8c",x"44",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"40",x"40",x"20",x"40",x"40",x"80",x"80",x"40",x"00",x"04",x"24",x"a4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"40",x"60",x"a0",x"c9",x"f2",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f6",x"cd",x"64",x"40",x"40",x"64",x"ad",x"cd",x"ed",x"ed",x"e9",x"e9",x"e9",x"e4",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"64",x"64",x"84",x"84",x"84",x"84",x"a5",x"a9",x"a9",x"cd",x"cd",x"cd",x"ed",x"ed",x"e9",x"c9",x"c5",x"a4",x"60",x"60",x"40",x"40",x"40",x"40",x"60",x"80",x"80",x"80",x"80",x"60",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"8c",x"d4",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f4",x"d0",x"b0",x"8c",x"a8",x"a4",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c8",x"f0",x"f8",x"fc",x"fc",x"fc",x"fd",x"fd",x"fe",x"ff",x"ff",x"ff",x"fe",x"fd",x"fc",x"fc",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"d0",x"d0",x"b0",x"b0",x"ac",x"8c",x"8c",x"8c",x"6c",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"d0",x"d4",x"d5",x"f5",x"f9",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"f8",x"f8",x"d4",x"d4",x"d0",x"cc",x"c8",x"a8",x"a4",x"c0",x"a0",x"80",x"80",x"80",x"80",x"64",x"a8",x"d0",x"b0",x"b0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d0",x"b0",x"b0",x"b0",x"ac",x"8c",x"84",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"c0",x"a0",x"c0",x"e0",x"c0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"c0",x"e0",x"c0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"64",x"88",x"ac",x"d0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"b0",x"ac",x"84",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"44",x"64",x"68",x"88",x"88",x"8c",x"8c",x"8c",x"ac",x"b0",x"d0",x"d4",x"d4",x"f4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"f9",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"d4",x"d4",x"d4",x"d0",x"d0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f9",x"f9",x"fd",x"fd",x"f9",x"f9",x"d4",x"d4",x"d4",x"d4",x"b0",x"b0",x"8c",x"64",x"40",x"40",x"40",x"40",x"40",x"20",x"44",x"68",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"b4",x"d4",x"d4",x"f8",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"f9",x"f9",x"f8",x"f8",x"f8",x"d4",x"d4",x"d4",x"d4",x"8c",x"64",x"40",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"40",x"40",x"40",x"20",x"40",x"60",x"80",x"60",x"20",x"04",x"24",x"64",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"80",x"a0",x"cd",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"a9",x"84",x"40",x"40",x"60",x"a9",x"cd",x"ed",x"ed",x"e9",x"e9",x"e4",x"e4",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"84",x"84",x"a4",x"a9",x"a9",x"c9",x"c9",x"cd",x"ed",x"ed",x"c9",x"c9",x"c9",x"a4",x"a4",x"80",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"80",x"80",x"60",x"60",x"40",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"40",x"60",x"88",x"d4",x"f9",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"d4",x"b4",x"b0",x"a8",x"a4",x"c4",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c4",x"ec",x"f4",x"f8",x"fc",x"fc",x"fd",x"fd",x"fd",x"fe",x"ff",x"ff",x"fe",x"fe",x"fd",x"fc",x"fc",x"f8",x"f8",x"f4",x"f5",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"b0",x"b0",x"8c",x"8c",x"8c",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"48",x"68",x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"68",x"6c",x"6c",x"6c",x"8c",x"8c",x"90",x"b0",x"b0",x"b0",x"d0",x"d4",x"d5",x"f5",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"fd",x"fd",x"f9",x"f8",x"d4",x"d4",x"d0",x"d0",x"ac",x"a8",x"a4",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"64",x"a8",x"cc",x"b0",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d0",x"d0",x"b0",x"b0",x"ac",x"8c",x"84",x"80",x"80",x"80",x"a0",x"c0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"c0",x"a0",x"c0",x"e0",x"c0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"c0",x"c0",x"c0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"64",x"88",x"ac",x"d0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"b0",x"ac",x"84",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"44",x"64",x"68",x"88",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"d5",x"d4",x"b0",x"b0",x"b0",x"b0",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"f9",x"f9",x"d4",x"d4",x"d4",x"d0",x"b0",x"b0",x"88",x"64",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"68",x"68",x"8c",x"8c",x"8c",x"90",x"b0",x"b0",x"b4",x"d4",x"d4",x"f8",x"f9",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fe",x"f9",x"f8",x"f8",x"f8",x"d4",x"d4",x"d4",x"d4",x"8c",x"68",x"40",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"60",x"80",x"80",x"40",x"20",x"04",x"44",x"84",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"80",x"60",x"40",x"60",x"60",x"80",x"a5",x"f2",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"d6",x"89",x"40",x"40",x"60",x"84",x"c9",x"e9",x"e9",x"e9",x"e5",x"e5",x"e4",x"e4",x"e4",x"c0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"84",x"a5",x"a5",x"a9",x"a9",x"cd",x"cd",x"ed",x"ed",x"e9",x"e9",x"e5",x"c4",x"80",x"60",x"60",x"40",x"20",x"40",x"40",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"60",x"60",x"60",x"40",x"40",x"40",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"64",x"88",x"d0",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"d8",x"d4",x"d4",x"b0",x"ac",x"c8",x"c4",x"c4",x"c0",x"c0",x"e0",x"e0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e8",x"f4",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fe",x"fe",x"ff",x"fe",x"fe",x"fe",x"fd",x"fc",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"b0",x"ac",x"8c",x"8c",x"8c",x"68",x"68",x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"44",x"44",x"44",x"44",x"44",x"48",x"48",x"68",x"68",x"68",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"d0",x"d5",x"f5",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"f9",x"f8",x"f4",x"f4",x"d4",x"d4",x"d0",x"ac",x"a4",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"a8",x"ac",x"b0",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"b0",x"b0",x"b0",x"ac",x"a8",x"84",x"80",x"80",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"64",x"88",x"ac",x"d0",x"d0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f5",x"d4",x"d0",x"b0",x"b0",x"b0",x"ac",x"84",x"80",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"64",x"68",x"88",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"f9",x"f9",x"f9",x"d4",x"b0",x"b0",x"b0",x"b0",x"b0",x"d0",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"f9",x"fd",x"fd",x"f9",x"f9",x"d4",x"d4",x"b0",x"b0",x"b0",x"8c",x"88",x"60",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"64",x"68",x"8c",x"8c",x"8c",x"90",x"b0",x"b0",x"b4",x"d4",x"d4",x"f8",x"f9",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fe",x"f9",x"f8",x"f8",x"f8",x"f8",x"d4",x"d4",x"d4",x"b0",x"68",x"44",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"80",x"a0",x"60",x"20",x"04",x"04",x"64",x"a4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"84",x"80",x"80",x"80",x"80",x"60",x"40",x"60",x"80",x"a0",x"a9",x"f6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d2",x"69",x"44",x"40",x"60",x"a4",x"c9",x"e9",x"e9",x"e9",x"e5",x"e4",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"84",x"84",x"84",x"85",x"a9",x"c9",x"e9",x"c9",x"c9",x"c9",x"c9",x"c9",x"c9",x"c4",x"a4",x"a0",x"80",x"60",x"60",x"40",x"40",x"20",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"88",x"d0",x"f8",x"f8",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"f9",x"f8",x"d8",x"d4",x"d4",x"d0",x"ac",x"ac",x"a8",x"c4",x"c0",x"e0",x"c0",x"c0",x"e0",x"e0",x"c0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"e0",x"e0",x"c0",x"e8",x"f0",x"f8",x"fc",x"fc",x"fc",x"fc",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d0",x"d0",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"6c",x"68",x"68",x"48",x"48",x"48",x"48",x"48",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"64",x"64",x"64",x"68",x"68",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"f9",x"f8",x"f4",x"f4",x"d4",x"d4",x"d0",x"cc",x"a8",x"a4",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"88",x"ac",x"b0",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"b0",x"b0",x"b0",x"ac",x"ac",x"88",x"84",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"c0",x"c0",x"c0",x"a0",x"c0",x"c0",x"a0",x"a0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"64",x"88",x"b0",x"d4",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"b0",x"ac",x"84",x"80",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"44",x"64",x"68",x"68",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"d0",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"d4",x"b0",x"b0",x"b0",x"8c",x"b0",x"b0",x"b0",x"d0",x"d4",x"d4",x"d4",x"d4",x"d4",x"f5",x"f9",x"f9",x"f9",x"d4",x"d4",x"b0",x"b0",x"b0",x"8c",x"8c",x"68",x"60",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"44",x"68",x"8c",x"8c",x"8c",x"90",x"90",x"b0",x"b0",x"b4",x"d4",x"d4",x"f9",x"f9",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fe",x"f9",x"f8",x"f8",x"f8",x"d4",x"d4",x"d4",x"d4",x"b0",x"8c",x"44",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"80",x"a0",x"60",x"04",x"04",x"24",x"84",x"c4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"80",x"80",x"80",x"60",x"80",x"80",x"60",x"40",x"60",x"a0",x"a5",x"b2",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"cd",x"84",x"20",x"40",x"80",x"c4",x"e9",x"e9",x"e9",x"e5",x"e4",x"e4",x"e4",x"e0",x"c0",x"a0",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"84",x"a8",x"a9",x"a9",x"cd",x"cd",x"ed",x"ed",x"e9",x"e9",x"c9",x"a4",x"80",x"60",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"84",x"ac",x"d4",x"fc",x"f8",x"fc",x"fc",x"fd",x"fe",x"fe",x"fe",x"fd",x"fc",x"fc",x"fc",x"fd",x"fd",x"fe",x"fe",x"fd",x"f8",x"d8",x"d4",x"d0",x"d0",x"b0",x"b0",x"8c",x"a8",x"c0",x"e0",x"c0",x"c0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c4",x"ec",x"f8",x"f8",x"fc",x"fc",x"fc",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"d0",x"d0",x"b0",x"ac",x"8c",x"8c",x"8c",x"8c",x"68",x"68",x"68",x"48",x"48",x"48",x"48",x"44",x"44",x"64",x"64",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"64",x"64",x"68",x"88",x"88",x"8c",x"8c",x"90",x"b0",x"b0",x"b0",x"d0",x"d4",x"f4",x"f4",x"f5",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d0",x"d0",x"b0",x"ac",x"a8",x"a4",x"a0",x"a0",x"80",x"80",x"60",x"64",x"88",x"ac",x"d0",x"b0",x"b0",x"d0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"ac",x"b0",x"ac",x"a8",x"a4",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"c0",x"c0",x"c0",x"a0",x"c0",x"a0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"84",x"a8",x"b0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f4",x"f4",x"d4",x"b0",x"b0",x"b0",x"b0",x"ac",x"84",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"64",x"64",x"68",x"68",x"8c",x"8c",x"8c",x"8c",x"ac",x"ac",x"b0",x"b0",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"ff",x"ff",x"ff",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"fd",x"f9",x"f9",x"f9",x"d5",x"d0",x"b0",x"ac",x"8c",x"8c",x"8c",x"8c",x"ac",x"b0",x"b0",x"d0",x"d0",x"d0",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"b0",x"b0",x"b0",x"b0",x"8c",x"88",x"68",x"64",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"64",x"8c",x"8c",x"8c",x"90",x"90",x"b0",x"b0",x"b0",x"d4",x"d4",x"f8",x"f9",x"f9",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fa",x"f9",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"b0",x"64",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"40",x"20",x"40",x"40",x"20",x"20",x"40",x"80",x"80",x"80",x"40",x"04",x"24",x"64",x"c4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"80",x"80",x"80",x"64",x"64",x"60",x"60",x"60",x"80",x"a0",x"cd",x"da",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"f7",x"ce",x"84",x"60",x"60",x"80",x"c4",x"e4",x"e5",x"e5",x"e4",x"e4",x"e4",x"e0",x"c0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"80",x"80",x"84",x"84",x"84",x"84",x"a9",x"a9",x"c9",x"cd",x"ed",x"ed",x"e9",x"c9",x"c9",x"a5",x"a4",x"84",x"80",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"80",x"80",x"80",x"88",x"b0",x"f8",x"fc",x"fc",x"fc",x"fc",x"fd",x"fe",x"fe",x"fe",x"fd",x"fc",x"fc",x"fc",x"fd",x"fd",x"fe",x"fe",x"fd",x"f8",x"d8",x"d4",x"d0",x"d0",x"b0",x"b0",x"8c",x"a8",x"c4",x"e0",x"c0",x"c0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c8",x"f0",x"f8",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fc",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"d0",x"b0",x"b0",x"8c",x"8c",x"8c",x"6c",x"68",x"68",x"68",x"48",x"48",x"48",x"44",x"44",x"44",x"64",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"64",x"64",x"68",x"88",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"b0",x"d0",x"d4",x"f4",x"f5",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"d0",x"d0",x"b0",x"ac",x"a4",x"a0",x"a0",x"a0",x"80",x"60",x"64",x"88",x"ac",x"d0",x"b0",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"ac",x"b0",x"ac",x"a8",x"a4",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"60",x"84",x"ac",x"b0",x"d4",x"f4",x"f4",x"f8",x"f8",x"fd",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f4",x"f4",x"d4",x"b0",x"b0",x"b0",x"ac",x"a8",x"84",x"60",x"80",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"64",x"68",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"ac",x"b0",x"b0",x"d0",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"d5",x"d0",x"b0",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"d0",x"d0",x"d0",x"b0",x"b0",x"b0",x"90",x"90",x"8c",x"8c",x"68",x"64",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"44",x"88",x"8c",x"8c",x"90",x"90",x"90",x"b0",x"b0",x"d4",x"d4",x"f8",x"f9",x"f9",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fa",x"f9",x"d8",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"b0",x"68",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"20",x"60",x"80",x"60",x"40",x"20",x"04",x"44",x"84",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"80",x"80",x"80",x"80",x"64",x"64",x"40",x"60",x"80",x"a0",x"a5",x"d2",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"cd",x"84",x"20",x"40",x"a4",x"e5",x"e9",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"80",x"80",x"80",x"80",x"60",x"64",x"85",x"a9",x"a9",x"a9",x"c9",x"cd",x"ed",x"ed",x"e9",x"e9",x"c4",x"a4",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"a8",x"d0",x"f8",x"fc",x"fc",x"fc",x"fc",x"fd",x"fe",x"fe",x"fe",x"fd",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"f9",x"f8",x"d4",x"d4",x"d0",x"b0",x"b0",x"b0",x"ac",x"a8",x"a4",x"c0",x"e0",x"e0",x"c0",x"c0",x"e0",x"c0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"c4",x"ec",x"f0",x"f8",x"f8",x"fc",x"fc",x"fc",x"fd",x"fd",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"d0",x"b0",x"b0",x"ac",x"8c",x"8c",x"68",x"68",x"68",x"48",x"48",x"48",x"44",x"44",x"44",x"44",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"64",x"64",x"68",x"88",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"d0",x"d0",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"ac",x"a8",x"a0",x"a0",x"a0",x"80",x"60",x"60",x"84",x"ac",x"d0",x"b0",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"b0",x"b0",x"b0",x"ac",x"a8",x"a4",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"c0",x"e0",x"c0",x"a0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"a0",x"c0",x"a0",x"a0",x"c0",x"c0",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"88",x"ac",x"b0",x"d0",x"d4",x"f4",x"f8",x"f9",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"b0",x"b0",x"b0",x"ac",x"a8",x"64",x"60",x"80",x"60",x"60",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"64",x"48",x"68",x"88",x"8c",x"8c",x"8c",x"8c",x"ac",x"b0",x"b0",x"b0",x"d0",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"d9",x"d4",x"b0",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"90",x"90",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"8c",x"68",x"68",x"64",x"40",x"60",x"60",x"40",x"40",x"60",x"60",x"40",x"20",x"40",x"44",x"68",x"8c",x"8c",x"90",x"90",x"90",x"b0",x"b0",x"d4",x"d4",x"d4",x"f8",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fe",x"f9",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"b0",x"68",x"40",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"60",x"40",x"40",x"40",x"60",x"60",x"80",x"40",x"00",x"00",x"44",x"84",x"c5",x"e4",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"80",x"84",x"80",x"80",x"60",x"24",x"60",x"a0",x"c0",x"c9",x"f6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d2",x"64",x"40",x"40",x"80",x"e4",x"e5",x"e5",x"e4",x"e4",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"84",x"88",x"a9",x"a9",x"c9",x"c9",x"e9",x"e9",x"c9",x"c5",x"a4",x"84",x"80",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"a0",x"80",x"80",x"a8",x"f0",x"f8",x"fc",x"fc",x"fc",x"fc",x"fd",x"fe",x"fe",x"fe",x"fd",x"fd",x"fc",x"fc",x"fc",x"fd",x"fd",x"f9",x"f9",x"f8",x"d4",x"d4",x"d0",x"b0",x"b0",x"b0",x"8c",x"ac",x"a4",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"c0",x"c0",x"c0",x"a0",x"a0",x"c8",x"f0",x"f4",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"fd",x"fe",x"fe",x"fd",x"fd",x"fd",x"fc",x"f8",x"f8",x"f4",x"d4",x"d4",x"d0",x"b0",x"b0",x"ac",x"8c",x"8c",x"8c",x"68",x"68",x"48",x"48",x"44",x"44",x"44",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"64",x"64",x"88",x"8c",x"8c",x"8c",x"ac",x"b0",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d0",x"b0",x"b0",x"ac",x"a8",x"a4",x"a0",x"80",x"80",x"80",x"60",x"64",x"ac",x"d0",x"b0",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"ac",x"ac",x"a8",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"80",x"80",x"80",x"80",x"60",x"60",x"ac",x"d0",x"d0",x"d0",x"d4",x"f4",x"f9",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"b0",x"b0",x"b0",x"ac",x"88",x"84",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"64",x"68",x"88",x"8c",x"8c",x"8c",x"8c",x"8c",x"90",x"b0",x"b0",x"b0",x"d0",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"fd",x"fd",x"f9",x"f9",x"f9",x"d5",x"d4",x"b0",x"b0",x"90",x"8c",x"8c",x"6c",x"6c",x"6c",x"6c",x"8c",x"90",x"90",x"b0",x"b0",x"90",x"90",x"90",x"90",x"90",x"90",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"68",x"68",x"64",x"40",x"40",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"44",x"68",x"6c",x"8c",x"90",x"90",x"90",x"b0",x"b0",x"b0",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fe",x"fd",x"f9",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"b0",x"8c",x"44",x"20",x"00",x"20",x"20",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"40",x"60",x"40",x"20",x"60",x"80",x"80",x"60",x"20",x"00",x"20",x"64",x"a5",x"e5",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"80",x"80",x"84",x"84",x"80",x"60",x"40",x"40",x"60",x"c0",x"c5",x"d2",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"ee",x"a5",x"20",x"20",x"a0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"c0",x"a0",x"80",x"60",x"60",x"80",x"80",x"80",x"84",x"64",x"84",x"a9",x"a9",x"a9",x"c9",x"c9",x"e9",x"e9",x"c5",x"a1",x"80",x"40",x"40",x"20",x"40",x"40",x"60",x"80",x"80",x"60",x"60",x"40",x"40",x"40",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"cc",x"f4",x"f8",x"f8",x"fc",x"fc",x"fc",x"fd",x"fe",x"fe",x"fe",x"fd",x"fd",x"fc",x"fc",x"fc",x"f9",x"f9",x"f9",x"f8",x"f8",x"d4",x"d4",x"b0",x"b0",x"b0",x"b0",x"8c",x"8c",x"a8",x"a4",x"a0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"a0",x"a0",x"cc",x"f4",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f4",x"d4",x"d0",x"b0",x"b0",x"ac",x"8c",x"8c",x"8c",x"68",x"68",x"68",x"48",x"28",x"24",x"44",x"40",x"40",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"80",x"60",x"60",x"60",x"80",x"60",x"60",x"60",x"80",x"60",x"60",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"64",x"64",x"88",x"88",x"8c",x"ac",x"ac",x"b0",x"b0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d0",x"b0",x"b0",x"ac",x"ac",x"a4",x"80",x"80",x"80",x"80",x"60",x"64",x"a8",x"d0",x"b0",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"d0",x"b0",x"b0",x"ac",x"a8",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"c0",x"a0",x"80",x"a0",x"c0",x"c0",x"a0",x"a0",x"80",x"a0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"60",x"80",x"c0",x"a0",x"60",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"60",x"64",x"cc",x"d0",x"d0",x"d4",x"d4",x"f9",x"fd",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f8",x"f4",x"d4",x"d0",x"b0",x"b0",x"b0",x"ac",x"88",x"80",x"60",x"60",x"60",x"80",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"60",x"64",x"68",x"88",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"d0",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"d4",x"b4",x"b0",x"90",x"8c",x"8c",x"8c",x"6c",x"68",x"68",x"68",x"6c",x"8c",x"8c",x"90",x"90",x"90",x"90",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"68",x"68",x"64",x"44",x"40",x"40",x"40",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"68",x"8c",x"8c",x"90",x"90",x"b0",x"b0",x"b0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"f9",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"b0",x"8c",x"44",x"20",x"00",x"20",x"20",x"00",x"00",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"a0",x"80",x"40",x"00",x"00",x"44",x"a4",x"c5",x"e5",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"64",x"64",x"64",x"84",x"84",x"80",x"40",x"40",x"60",x"80",x"c0",x"c9",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"ce",x"85",x"60",x"60",x"80",x"c4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"60",x"60",x"80",x"80",x"80",x"84",x"88",x"88",x"cd",x"ed",x"e9",x"e9",x"c9",x"a4",x"84",x"80",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"c0",x"a0",x"a0",x"cc",x"f4",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fd",x"fe",x"fe",x"fd",x"fd",x"fc",x"fc",x"f8",x"f8",x"f9",x"f9",x"f8",x"f8",x"f4",x"d4",x"d0",x"b0",x"b0",x"b0",x"b0",x"8c",x"88",x"a4",x"c0",x"c0",x"c0",x"a0",x"c0",x"a0",x"80",x"a0",x"c0",x"c0",x"a0",x"a0",x"a4",x"cc",x"f8",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"8c",x"6c",x"68",x"68",x"48",x"44",x"44",x"44",x"40",x"40",x"60",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"64",x"64",x"88",x"88",x"8c",x"ac",x"b0",x"b0",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d0",x"b0",x"b0",x"b0",x"ac",x"a8",x"a4",x"80",x"80",x"80",x"60",x"60",x"88",x"ac",x"b0",x"b0",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"ac",x"a8",x"a4",x"a0",x"a0",x"a0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"88",x"d0",x"f4",x"d4",x"d4",x"d4",x"f9",x"fd",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f8",x"f8",x"f4",x"d4",x"b0",x"b0",x"b0",x"ac",x"ac",x"88",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"68",x"68",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"b0",x"d0",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"d5",x"d4",x"b0",x"b0",x"90",x"90",x"8c",x"8c",x"6c",x"68",x"68",x"48",x"48",x"68",x"68",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"68",x"68",x"44",x"44",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"44",x"68",x"8c",x"8c",x"90",x"90",x"b0",x"b0",x"b0",x"d4",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"f9",x"f9",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"b4",x"8c",x"48",x"20",x"00",x"00",x"00",x"00",x"00",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"60",x"80",x"80",x"60",x"20",x"00",x"24",x"64",x"c5",x"e5",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"64",x"64",x"84",x"84",x"84",x"60",x"40",x"60",x"a0",x"c0",x"c4",x"d2",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ee",x"a4",x"40",x"40",x"a4",x"e4",x"e5",x"e4",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"60",x"60",x"80",x"80",x"a0",x"a4",x"a4",x"a9",x"ad",x"ed",x"ed",x"e9",x"c5",x"a4",x"60",x"40",x"20",x"20",x"40",x"60",x"60",x"60",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"ec",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"fe",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"b0",x"b0",x"b0",x"b0",x"ac",x"68",x"84",x"c0",x"c0",x"a0",x"a0",x"c0",x"a0",x"80",x"a0",x"c0",x"c0",x"a0",x"a0",x"a8",x"d0",x"f8",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"f8",x"f8",x"f4",x"d4",x"d4",x"d0",x"d0",x"b0",x"8c",x"8c",x"6c",x"6c",x"6c",x"68",x"68",x"48",x"44",x"44",x"40",x"40",x"40",x"60",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"80",x"60",x"60",x"60",x"80",x"60",x"60",x"60",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"64",x"88",x"8c",x"ac",x"b0",x"b0",x"b0",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"b0",x"b0",x"90",x"b0",x"a8",x"a4",x"80",x"80",x"80",x"80",x"80",x"88",x"ac",x"b0",x"d0",x"b0",x"d0",x"d0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"d4",x"b4",x"b0",x"b0",x"ac",x"ac",x"88",x"84",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"c0",x"a0",x"60",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"a4",x"ac",x"d0",x"d4",x"f4",x"f4",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f8",x"f9",x"f4",x"d4",x"b0",x"b0",x"b0",x"ac",x"ac",x"88",x"60",x"60",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"64",x"68",x"68",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"b0",x"d0",x"d0",x"d0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"d4",x"d4",x"b0",x"b0",x"90",x"90",x"8c",x"8c",x"8c",x"8c",x"68",x"68",x"44",x"44",x"44",x"44",x"68",x"68",x"68",x"8c",x"8c",x"6c",x"6c",x"6c",x"6c",x"6c",x"8c",x"8c",x"8c",x"88",x"68",x"68",x"44",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"40",x"40",x"60",x"60",x"40",x"20",x"40",x"40",x"40",x"64",x"8c",x"8c",x"90",x"90",x"b0",x"b0",x"b0",x"b0",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"f9",x"f9",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"b4",x"90",x"68",x"24",x"00",x"00",x"00",x"00",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"a0",x"80",x"60",x"20",x"00",x"24",x"64",x"a9",x"e5",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"80",x"84",x"84",x"84",x"84",x"80",x"60",x"40",x"60",x"c0",x"c4",x"cd",x"d6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d2",x"85",x"60",x"40",x"80",x"c4",x"e4",x"e4",x"e0",x"e0",x"e0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"80",x"84",x"a4",x"a9",x"c9",x"cd",x"cd",x"e9",x"c8",x"a4",x"80",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e8",x"f0",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"fe",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"b0",x"b0",x"b0",x"b0",x"8c",x"8c",x"84",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"a0",x"c0",x"a0",x"a0",x"a4",x"cc",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"f8",x"f8",x"f4",x"d4",x"d4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"68",x"6c",x"68",x"68",x"44",x"44",x"44",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"84",x"88",x"ac",x"ac",x"b0",x"b0",x"b0",x"b0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"b0",x"b0",x"b0",x"b0",x"ac",x"a8",x"80",x"80",x"80",x"60",x"60",x"84",x"8c",x"ac",x"b0",x"b0",x"d0",x"d0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"b0",x"ac",x"a8",x"a4",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"a0",x"80",x"80",x"80",x"a8",x"cc",x"d4",x"d4",x"f4",x"f8",x"f9",x"fd",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f9",x"f9",x"f5",x"d4",x"b0",x"ac",x"ac",x"8c",x"88",x"84",x"60",x"60",x"60",x"60",x"80",x"60",x"60",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"48",x"68",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"90",x"b0",x"b0",x"b0",x"b0",x"d0",x"d0",x"d0",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"d4",x"d4",x"b0",x"b0",x"90",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"68",x"68",x"44",x"40",x"40",x"40",x"40",x"44",x"44",x"64",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"64",x"44",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"20",x"20",x"44",x"8c",x"8c",x"90",x"90",x"90",x"b0",x"b0",x"b0",x"d4",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"f9",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"b4",x"90",x"6c",x"24",x"00",x"00",x"00",x"20",x"40",x"20",x"20",x"40",x"60",x"40",x"40",x"40",x"60",x"80",x"60",x"20",x"00",x"00",x"64",x"a9",x"e9",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"80",x"84",x"84",x"84",x"64",x"60",x"60",x"80",x"a0",x"c0",x"c9",x"f6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"d2",x"a5",x"40",x"40",x"80",x"c0",x"e4",x"e4",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"85",x"a9",x"cd",x"ed",x"ed",x"c9",x"a4",x"80",x"40",x"40",x"20",x"20",x"40",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e8",x"f0",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"b0",x"b0",x"b0",x"90",x"8c",x"8c",x"88",x"80",x"a0",x"c0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"80",x"a8",x"d0",x"f8",x"f8",x"fc",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"d0",x"d0",x"b0",x"ac",x"8c",x"6c",x"68",x"68",x"68",x"48",x"44",x"64",x"60",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"64",x"84",x"a8",x"ac",x"b0",x"b0",x"b0",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"b4",x"b0",x"b0",x"b0",x"ac",x"88",x"84",x"a0",x"80",x"60",x"60",x"84",x"88",x"ac",x"b0",x"b0",x"d0",x"d0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"f4",x"f4",x"d4",x"b0",x"b0",x"b0",x"cc",x"a8",x"84",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"60",x"80",x"a0",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"a4",x"cc",x"d0",x"d4",x"d4",x"f4",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f9",x"f9",x"f5",x"d0",x"b0",x"ac",x"8c",x"8c",x"88",x"64",x"80",x"60",x"60",x"60",x"80",x"80",x"60",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"44",x"68",x"68",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"b0",x"d0",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"d4",x"d4",x"b4",x"b0",x"90",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"88",x"64",x"44",x"40",x"40",x"20",x"20",x"40",x"40",x"40",x"40",x"44",x"44",x"44",x"64",x"64",x"64",x"64",x"64",x"64",x"64",x"44",x"40",x"40",x"20",x"20",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"60",x"40",x"40",x"60",x"60",x"40",x"20",x"20",x"44",x"88",x"8c",x"90",x"90",x"90",x"b0",x"b0",x"b0",x"d4",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"f9",x"f5",x"f4",x"f4",x"f4",x"d4",x"d4",x"b4",x"90",x"6c",x"24",x"00",x"00",x"00",x"40",x"40",x"20",x"20",x"40",x"60",x"40",x"40",x"80",x"80",x"80",x"40",x"00",x"00",x"24",x"84",x"e9",x"e5",x"e4",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"84",x"84",x"84",x"60",x"40",x"60",x"a0",x"a0",x"a0",x"cd",x"fb",x"ff",x"ff",x"ff",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"f6",x"89",x"60",x"40",x"60",x"c0",x"e0",x"e4",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"80",x"84",x"84",x"84",x"85",x"c9",x"ed",x"ed",x"e9",x"c9",x"84",x"40",x"20",x"40",x"40",x"40",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"64",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"64",x"64",x"44",x"44",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c8",x"f0",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"d4",x"d4",x"b0",x"b0",x"b0",x"8c",x"8c",x"88",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"a0",x"a0",x"a0",x"80",x"c8",x"f4",x"f8",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"f8",x"f8",x"f8",x"f4",x"d4",x"d0",x"d0",x"b0",x"b0",x"8c",x"8c",x"68",x"68",x"68",x"68",x"44",x"44",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"64",x"88",x"ac",x"ac",x"b0",x"b0",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"b0",x"b0",x"b0",x"b0",x"a8",x"a4",x"80",x"80",x"80",x"60",x"60",x"84",x"ac",x"b0",x"b0",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"d0",x"d0",x"d0",x"ac",x"84",x"80",x"80",x"80",x"80",x"80",x"a0",x"80",x"80",x"80",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"a4",x"a8",x"d0",x"d4",x"d4",x"f4",x"f8",x"f9",x"fd",x"fd",x"fd",x"fd",x"f9",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f8",x"f9",x"f9",x"f4",x"d0",x"b0",x"8c",x"8c",x"8c",x"88",x"64",x"60",x"60",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"40",x"44",x"44",x"68",x"68",x"68",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f5",x"f5",x"f5",x"f5",x"d5",x"d4",x"d4",x"d4",x"b0",x"b0",x"b0",x"90",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"68",x"68",x"64",x"64",x"40",x"40",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"20",x"20",x"40",x"68",x"8c",x"8c",x"90",x"90",x"b0",x"b0",x"b0",x"b4",x"d4",x"d4",x"f8",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"f9",x"f9",x"f4",x"f8",x"f4",x"d4",x"d4",x"d4",x"b0",x"6c",x"24",x"00",x"20",x"40",x"40",x"40",x"20",x"20",x"20",x"40",x"60",x"80",x"a0",x"80",x"20",x"00",x"00",x"24",x"68",x"c9",x"e5",x"e4",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"80",x"a4",x"84",x"60",x"60",x"60",x"80",x"c0",x"c0",x"a9",x"d6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"f7",x"ce",x"64",x"40",x"60",x"a0",x"e4",x"e4",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"60",x"80",x"80",x"84",x"84",x"64",x"89",x"a9",x"ed",x"ed",x"e9",x"c9",x"80",x"40",x"00",x"00",x"40",x"60",x"60",x"80",x"60",x"60",x"40",x"40",x"40",x"44",x"64",x"48",x"68",x"6c",x"8c",x"b0",x"b0",x"b0",x"b4",x"b4",x"b4",x"b4",x"b4",x"b4",x"b4",x"d0",x"d0",x"d0",x"b0",x"b0",x"8c",x"8c",x"8c",x"88",x"68",x"64",x"64",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c4",x"cc",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"b0",x"b0",x"b0",x"b0",x"6c",x"68",x"a4",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a4",x"cc",x"f5",x"f8",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"d0",x"b0",x"ac",x"8c",x"8c",x"68",x"68",x"68",x"48",x"44",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"84",x"88",x"ac",x"ac",x"b0",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f0",x"d0",x"b0",x"b0",x"b0",x"ac",x"a8",x"80",x"60",x"80",x"80",x"60",x"64",x"8c",x"ac",x"ac",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"f4",x"f4",x"d0",x"d0",x"d0",x"b0",x"88",x"80",x"80",x"80",x"80",x"80",x"a0",x"80",x"80",x"80",x"a0",x"80",x"60",x"80",x"a0",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"a4",x"cc",x"d4",x"f4",x"f4",x"f4",x"f8",x"f9",x"fd",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f9",x"f9",x"f9",x"d4",x"b0",x"b0",x"8c",x"8c",x"88",x"84",x"60",x"60",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"40",x"44",x"64",x"68",x"68",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"d8",x"d8",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"b0",x"b0",x"b0",x"90",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"68",x"68",x"68",x"64",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"20",x"40",x"44",x"68",x"8c",x"8c",x"8c",x"90",x"b0",x"b0",x"b0",x"d4",x"d4",x"f4",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"fd",x"f9",x"f9",x"f4",x"f8",x"d4",x"d4",x"d4",x"b4",x"b0",x"6c",x"44",x"20",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"80",x"a0",x"a0",x"60",x"00",x"00",x"24",x"68",x"a9",x"e5",x"e4",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"84",x"84",x"a4",x"80",x"80",x"40",x"60",x"80",x"a0",x"c0",x"c5",x"b2",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"cd",x"a4",x"60",x"60",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"a0",x"a0",x"80",x"80",x"60",x"80",x"80",x"84",x"84",x"88",x"89",x"ad",x"ed",x"e9",x"e9",x"c4",x"80",x"40",x"20",x"40",x"40",x"40",x"40",x"40",x"60",x"64",x"88",x"8c",x"8c",x"b0",x"b0",x"b4",x"b4",x"d8",x"d8",x"d8",x"d8",x"d8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"d8",x"d8",x"d4",x"d4",x"d4",x"b0",x"b0",x"ac",x"a8",x"a8",x"a4",x"a4",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a4",x"a8",x"d0",x"f8",x"f4",x"f4",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"b0",x"b0",x"b0",x"ac",x"8c",x"88",x"84",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a8",x"d0",x"f5",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"8c",x"68",x"68",x"48",x"44",x"44",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"84",x"88",x"ac",x"b0",x"b0",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"b0",x"ac",x"a8",x"84",x"80",x"80",x"60",x"60",x"60",x"88",x"ac",x"ac",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"b0",x"ac",x"84",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"ac",x"d0",x"f4",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"fd",x"fd",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f8",x"f9",x"f9",x"f5",x"d0",x"b0",x"ac",x"8c",x"8c",x"88",x"64",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"64",x"68",x"88",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"90",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"b4",x"b0",x"b0",x"b0",x"b0",x"b0",x"90",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"68",x"68",x"64",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"44",x"68",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"d4",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"d4",x"d4",x"d4",x"d4",x"d4",x"b0",x"90",x"68",x"44",x"20",x"40",x"40",x"40",x"20",x"40",x"20",x"20",x"40",x"a0",x"a0",x"40",x"20",x"00",x"24",x"69",x"a9",x"e9",x"e5",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"80",x"84",x"84",x"84",x"a4",x"84",x"60",x"60",x"80",x"c0",x"c0",x"a4",x"cd",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d2",x"84",x"60",x"80",x"a0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"64",x"64",x"89",x"a9",x"ed",x"ed",x"e9",x"c0",x"80",x"40",x"20",x"40",x"60",x"80",x"60",x"40",x"44",x"68",x"8c",x"b0",x"d4",x"d8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f4",x"d0",x"d0",x"cc",x"c8",x"a4",x"a4",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a4",x"a8",x"d0",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f8",x"f4",x"d4",x"d4",x"b0",x"b0",x"b0",x"8c",x"ac",x"ac",x"84",x"80",x"a0",x"a0",x"80",x"a0",x"c0",x"a0",x"a0",x"a4",x"a8",x"d0",x"f5",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"d0",x"b0",x"ac",x"8c",x"8c",x"68",x"68",x"68",x"48",x"44",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"64",x"88",x"ac",x"ac",x"b0",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"d0",x"ac",x"8c",x"8c",x"8c",x"84",x"80",x"60",x"60",x"60",x"60",x"88",x"8c",x"ac",x"b0",x"d0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"ac",x"a4",x"a0",x"a0",x"80",x"80",x"80",x"a0",x"80",x"80",x"80",x"a0",x"80",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"a0",x"a0",x"60",x"60",x"a0",x"a0",x"60",x"60",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"ac",x"d0",x"f4",x"f4",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"f9",x"f8",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f5",x"f5",x"d0",x"b0",x"ac",x"8c",x"8c",x"68",x"64",x"60",x"80",x"80",x"60",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"64",x"68",x"68",x"68",x"68",x"6c",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"90",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"90",x"8c",x"8c",x"8c",x"8c",x"6c",x"6c",x"6c",x"8c",x"8c",x"68",x"68",x"68",x"64",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"48",x"8c",x"8c",x"8c",x"8c",x"90",x"b0",x"b0",x"b0",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"d5",x"d4",x"d4",x"d4",x"d4",x"b4",x"b0",x"8c",x"68",x"40",x"20",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"60",x"a0",x"80",x"20",x"00",x"04",x"44",x"a9",x"e9",x"e5",x"e4",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"84",x"84",x"84",x"84",x"84",x"64",x"60",x"60",x"a0",x"c0",x"c0",x"a9",x"d6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"b2",x"64",x"40",x"40",x"80",x"c0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"a0",x"80",x"64",x"68",x"68",x"a9",x"e9",x"e9",x"e5",x"a0",x"60",x"20",x"20",x"40",x"60",x"64",x"68",x"8c",x"b0",x"b4",x"d4",x"d8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f4",x"f4",x"d0",x"d0",x"cc",x"cc",x"c4",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"80",x"84",x"d0",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f8",x"f4",x"d4",x"d0",x"b0",x"b0",x"b0",x"ac",x"ac",x"ac",x"88",x"84",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"80",x"a4",x"cc",x"f0",x"f4",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"d0",x"b0",x"8c",x"8c",x"8c",x"68",x"68",x"68",x"44",x"44",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"84",x"88",x"ac",x"b0",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"f0",x"d0",x"d0",x"ac",x"8c",x"8c",x"8c",x"84",x"80",x"80",x"60",x"60",x"60",x"88",x"8c",x"ac",x"ac",x"b0",x"d0",x"d0",x"d0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"b4",x"d0",x"cc",x"a8",x"a0",x"80",x"80",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"80",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"a8",x"d0",x"f4",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"f9",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f5",x"d5",x"b0",x"ac",x"8c",x"8c",x"8c",x"68",x"64",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"44",x"68",x"68",x"68",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"ac",x"ac",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"6c",x"68",x"68",x"64",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"44",x"6c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f8",x"f9",x"f9",x"d5",x"d4",x"d4",x"b4",x"b4",x"b0",x"b0",x"8c",x"68",x"40",x"20",x"40",x"40",x"20",x"20",x"40",x"60",x"a0",x"a0",x"60",x"20",x"04",x"04",x"48",x"a9",x"e9",x"e9",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"80",x"80",x"84",x"a4",x"84",x"64",x"44",x"64",x"a0",x"c0",x"a0",x"c4",x"d2",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"89",x"40",x"40",x"60",x"a0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"84",x"48",x"69",x"8d",x"c9",x"e5",x"e4",x"c0",x"60",x"20",x"20",x"20",x"60",x"84",x"8c",x"90",x"b4",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f4",x"f4",x"f0",x"c8",x"c4",x"c4",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"84",x"ac",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f9",x"f8",x"f4",x"d4",x"d4",x"b0",x"b0",x"b0",x"ac",x"ac",x"8c",x"88",x"84",x"a0",x"a0",x"a0",x"a0",x"c0",x"a0",x"80",x"a4",x"d0",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"8c",x"68",x"68",x"48",x"44",x"44",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"60",x"64",x"88",x"ac",x"ac",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"f0",x"f0",x"d0",x"ac",x"8c",x"ac",x"ac",x"88",x"84",x"60",x"60",x"60",x"60",x"64",x"88",x"8c",x"ac",x"b0",x"d0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"d0",x"cc",x"a8",x"a0",x"80",x"a0",x"80",x"80",x"80",x"a0",x"80",x"80",x"80",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"a0",x"80",x"60",x"60",x"80",x"80",x"80",x"60",x"60",x"80",x"a0",x"80",x"84",x"cc",x"f5",x"f8",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"f9",x"f8",x"f8",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f5",x"d0",x"b0",x"ac",x"8c",x"8c",x"88",x"68",x"60",x"40",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"44",x"64",x"68",x"68",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"68",x"68",x"64",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"44",x"68",x"8c",x"8c",x"8c",x"8c",x"90",x"b0",x"b0",x"d4",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"d4",x"f9",x"f5",x"d4",x"d4",x"b4",x"b4",x"b0",x"b0",x"8c",x"88",x"64",x"40",x"20",x"40",x"40",x"20",x"20",x"40",x"80",x"c0",x"a0",x"20",x"00",x"04",x"48",x"a9",x"c9",x"e9",x"e5",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"a4",x"85",x"64",x"64",x"44",x"64",x"c0",x"c0",x"a0",x"a9",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"b2",x"64",x"20",x"60",x"a0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"80",x"80",x"60",x"80",x"80",x"80",x"84",x"65",x"69",x"8d",x"c9",x"e9",x"e4",x"a0",x"60",x"40",x"20",x"40",x"68",x"ac",x"d4",x"d8",x"d8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d0",x"cc",x"cc",x"c4",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"60",x"60",x"a8",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d0",x"b0",x"b0",x"b0",x"90",x"8c",x"88",x"84",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a8",x"d0",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"8c",x"8c",x"8c",x"8c",x"68",x"68",x"48",x"44",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"84",x"a8",x"ac",x"b0",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"d0",x"b0",x"ac",x"ac",x"ac",x"88",x"84",x"60",x"60",x"40",x"40",x"40",x"64",x"8c",x"ac",x"ac",x"b0",x"d0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"f4",x"f4",x"d4",x"d0",x"c8",x"a4",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"a4",x"a8",x"cc",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f8",x"f9",x"f9",x"f9",x"d5",x"b0",x"b0",x"8c",x"8c",x"88",x"88",x"64",x"40",x"40",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"64",x"64",x"64",x"68",x"68",x"68",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"88",x"68",x"68",x"64",x"64",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"44",x"68",x"8c",x"8c",x"8c",x"8c",x"90",x"b0",x"b0",x"b4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d0",x"d0",x"b0",x"b0",x"b0",x"90",x"8c",x"8c",x"68",x"44",x"40",x"40",x"20",x"20",x"40",x"60",x"80",x"80",x"60",x"20",x"00",x"04",x"49",x"8d",x"cd",x"e9",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a4",x"84",x"a4",x"a5",x"85",x"65",x"44",x"44",x"80",x"a0",x"a0",x"a0",x"c9",x"f2",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"d6",x"89",x"40",x"20",x"80",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"64",x"64",x"69",x"89",x"c9",x"e9",x"e4",x"c0",x"80",x"40",x"40",x"44",x"88",x"b0",x"d8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"d8",x"d4",x"d0",x"cc",x"a8",x"a4",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"88",x"b0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"d0",x"b0",x"b0",x"b0",x"90",x"90",x"6c",x"88",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c8",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"6c",x"48",x"44",x"44",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"80",x"80",x"60",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"84",x"a8",x"ac",x"b0",x"b0",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"b0",x"b0",x"8c",x"88",x"60",x"40",x"40",x"40",x"40",x"64",x"88",x"ac",x"ac",x"b0",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"cc",x"a8",x"84",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"64",x"84",x"ac",x"d0",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"fd",x"fd",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f8",x"f9",x"f9",x"d5",x"d0",x"b0",x"90",x"8c",x"8c",x"68",x"64",x"60",x"40",x"40",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"64",x"64",x"64",x"68",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"8c",x"6c",x"68",x"68",x"68",x"64",x"64",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"44",x"8c",x"8c",x"8c",x"8c",x"90",x"90",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"d0",x"d0",x"b4",x"b4",x"b4",x"b0",x"b0",x"ac",x"b0",x"b0",x"90",x"90",x"6c",x"68",x"44",x"40",x"40",x"40",x"20",x"40",x"60",x"80",x"80",x"60",x"20",x"00",x"04",x"49",x"8d",x"cd",x"e9",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"84",x"84",x"a4",x"a5",x"85",x"64",x"44",x"60",x"c0",x"c0",x"80",x"a4",x"f2",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"f6",x"8d",x"44",x"40",x"60",x"a0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"a0",x"80",x"44",x"44",x"64",x"a9",x"e9",x"e8",x"e4",x"a0",x"60",x"40",x"40",x"88",x"b0",x"d4",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d0",x"cc",x"a8",x"a8",x"a4",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"60",x"60",x"84",x"ac",x"d4",x"f8",x"f4",x"f8",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"b0",x"b0",x"ac",x"90",x"90",x"6c",x"68",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c8",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"b0",x"b0",x"8c",x"8c",x"8c",x"88",x"68",x"48",x"44",x"44",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"60",x"80",x"80",x"a0",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"64",x"a8",x"ac",x"b0",x"b0",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"b0",x"b0",x"ac",x"88",x"60",x"40",x"40",x"40",x"40",x"60",x"88",x"8c",x"ac",x"b0",x"b0",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"f4",x"f4",x"f0",x"cc",x"a8",x"84",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"60",x"60",x"60",x"80",x"a8",x"cc",x"d0",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"fd",x"fd",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f8",x"f8",x"f9",x"f5",x"d5",x"b0",x"b0",x"8c",x"8c",x"8c",x"88",x"44",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"64",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"88",x"8c",x"6c",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"6c",x"6c",x"6c",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"64",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"44",x"8c",x"8c",x"8c",x"8c",x"8c",x"90",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b4",x"b0",x"b0",x"ac",x"8c",x"ac",x"ac",x"8c",x"8c",x"6c",x"48",x"44",x"40",x"40",x"40",x"40",x"60",x"80",x"80",x"40",x"20",x"00",x"04",x"69",x"ad",x"cd",x"e9",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"64",x"64",x"84",x"85",x"85",x"64",x"44",x"60",x"80",x"c0",x"c0",x"a4",x"cd",x"f6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"ee",x"64",x"20",x"60",x"a0",x"c0",x"e0",x"e0",x"e0",x"c0",x"80",x"60",x"60",x"80",x"80",x"a0",x"84",x"44",x"48",x"89",x"c9",x"e4",x"e4",x"c0",x"80",x"40",x"64",x"88",x"d0",x"f8",x"fc",x"fc",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fe",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d0",x"d0",x"ac",x"a8",x"a4",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"64",x"88",x"d0",x"f8",x"f4",x"f4",x"f8",x"f8",x"f8",x"fc",x"fc",x"fd",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"b0",x"b0",x"ac",x"90",x"8c",x"6c",x"68",x"84",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c8",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"b0",x"b0",x"8c",x"8c",x"88",x"88",x"68",x"48",x"44",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"60",x"84",x"ac",x"b0",x"b0",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"b0",x"b0",x"ac",x"88",x"64",x"40",x"40",x"40",x"40",x"40",x"64",x"88",x"ac",x"b0",x"b0",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"f4",x"f4",x"f4",x"f4",x"d0",x"a8",x"84",x"80",x"60",x"60",x"60",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"80",x"80",x"64",x"84",x"84",x"a8",x"d0",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f8",x"f9",x"f9",x"d4",x"d4",x"b0",x"90",x"8c",x"8c",x"88",x"64",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"60",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"44",x"44",x"44",x"64",x"44",x"64",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"64",x"64",x"64",x"64",x"64",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"44",x"68",x"68",x"68",x"6c",x"8c",x"8c",x"90",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"90",x"90",x"8c",x"8c",x"8c",x"8c",x"ac",x"8c",x"8c",x"48",x"28",x"24",x"40",x"40",x"60",x"60",x"80",x"80",x"60",x"20",x"00",x"04",x"49",x"ad",x"d1",x"ed",x"e9",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"64",x"44",x"84",x"85",x"85",x"64",x"44",x"64",x"a0",x"c0",x"c0",x"c0",x"cd",x"d6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"f6",x"a5",x"60",x"20",x"80",x"c0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"60",x"80",x"80",x"84",x"64",x"48",x"88",x"cd",x"e8",x"e0",x"e0",x"a0",x"64",x"68",x"90",x"d8",x"f9",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fe",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f5",x"d0",x"b0",x"8c",x"84",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"68",x"d0",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"b0",x"b0",x"ac",x"8c",x"8c",x"8c",x"68",x"64",x"80",x"c0",x"a0",x"80",x"80",x"a0",x"c8",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"b0",x"b0",x"8c",x"8c",x"88",x"88",x"68",x"48",x"44",x"40",x"60",x"60",x"60",x"80",x"80",x"60",x"60",x"80",x"80",x"a0",x"80",x"80",x"80",x"a0",x"a0",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"c0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"60",x"60",x"64",x"88",x"b0",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"b0",x"ac",x"88",x"64",x"40",x"40",x"40",x"40",x"40",x"40",x"64",x"8c",x"ac",x"b0",x"b0",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f8",x"f8",x"f4",x"d4",x"d4",x"f4",x"f4",x"f4",x"d0",x"cc",x"a8",x"84",x"80",x"60",x"60",x"60",x"60",x"80",x"60",x"60",x"60",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"84",x"a8",x"cc",x"f1",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"fd",x"fd",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f9",x"f9",x"d5",x"d4",x"b0",x"b0",x"8c",x"8c",x"8c",x"68",x"44",x"60",x"60",x"40",x"40",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"60",x"40",x"60",x"80",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"40",x"44",x"44",x"64",x"64",x"44",x"64",x"64",x"64",x"64",x"64",x"64",x"64",x"44",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"44",x"44",x"68",x"68",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"b0",x"b0",x"90",x"70",x"70",x"8c",x"90",x"91",x"8c",x"68",x"44",x"20",x"20",x"20",x"60",x"80",x"80",x"80",x"40",x"20",x"20",x"44",x"6d",x"91",x"d1",x"ed",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"84",x"84",x"84",x"84",x"85",x"69",x"44",x"60",x"80",x"c0",x"e0",x"c0",x"a4",x"f6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"cd",x"80",x"40",x"40",x"a0",x"e0",x"e0",x"e0",x"e0",x"c0",x"80",x"60",x"60",x"60",x"80",x"80",x"64",x"69",x"89",x"a9",x"e8",x"e4",x"e0",x"c0",x"a0",x"88",x"94",x"d8",x"fc",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fe",x"fe",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"fc",x"f8",x"f9",x"f9",x"f4",x"d4",x"b0",x"88",x"84",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"80",x"60",x"60",x"60",x"40",x"64",x"b0",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"b0",x"b0",x"ac",x"ac",x"8c",x"8c",x"68",x"64",x"84",x"a0",x"a0",x"a0",x"a0",x"a0",x"c8",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"b0",x"b0",x"8c",x"8c",x"88",x"88",x"68",x"48",x"44",x"40",x"60",x"60",x"60",x"80",x"80",x"60",x"60",x"80",x"a0",x"a0",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"a0",x"c0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"40",x"40",x"40",x"40",x"64",x"88",x"b0",x"b0",x"d0",x"d0",x"d0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"b0",x"ac",x"88",x"64",x"60",x"40",x"40",x"40",x"40",x"40",x"64",x"88",x"ac",x"ac",x"b0",x"b0",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f8",x"d4",x"d4",x"f8",x"f8",x"f8",x"f4",x"f4",x"d0",x"ac",x"a8",x"84",x"84",x"80",x"84",x"84",x"64",x"60",x"80",x"80",x"84",x"84",x"80",x"80",x"84",x"84",x"88",x"a8",x"ec",x"f0",x"f5",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fd",x"fd",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f9",x"f5",x"d4",x"b0",x"90",x"90",x"8c",x"8c",x"88",x"44",x"40",x"60",x"60",x"40",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"80",x"60",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"44",x"48",x"68",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"6c",x"8c",x"8c",x"8c",x"68",x"64",x"40",x"40",x"40",x"40",x"80",x"80",x"80",x"60",x"20",x"20",x"49",x"6d",x"b2",x"d2",x"ed",x"e8",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"84",x"84",x"a8",x"a5",x"85",x"64",x"64",x"64",x"80",x"a0",x"c0",x"c0",x"c4",x"cd",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d2",x"89",x"40",x"60",x"80",x"c0",x"e0",x"e0",x"e0",x"c0",x"80",x"80",x"60",x"60",x"80",x"80",x"84",x"48",x"69",x"c5",x"e5",x"e0",x"c0",x"a0",x"a4",x"ac",x"d4",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fc",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d0",x"ac",x"a8",x"84",x"64",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"ac",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"b0",x"b0",x"ac",x"ac",x"8c",x"6c",x"6c",x"84",x"84",x"80",x"a0",x"a0",x"a0",x"84",x"ac",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"b0",x"b0",x"8c",x"8c",x"88",x"88",x"68",x"48",x"44",x"40",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"80",x"80",x"c0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"60",x"88",x"ac",x"b0",x"d0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"d0",x"b0",x"ac",x"ac",x"ac",x"84",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"88",x"8c",x"ac",x"b0",x"b0",x"b0",x"b0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"f8",x"f8",x"f4",x"f4",x"f4",x"f8",x"f8",x"f4",x"f4",x"d0",x"cc",x"ac",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"a8",x"cc",x"cc",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f9",x"f9",x"d5",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"68",x"64",x"60",x"40",x"40",x"60",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"24",x"44",x"48",x"68",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"48",x"44",x"40",x"40",x"40",x"40",x"60",x"80",x"a0",x"80",x"40",x"20",x"44",x"69",x"91",x"b2",x"ee",x"e9",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"80",x"64",x"64",x"89",x"a9",x"a5",x"84",x"64",x"64",x"64",x"c0",x"e0",x"c0",x"a0",x"ce",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"f6",x"a9",x"60",x"40",x"80",x"c0",x"e0",x"e0",x"e0",x"e0",x"a0",x"80",x"80",x"60",x"80",x"80",x"84",x"85",x"49",x"89",x"e5",x"e0",x"e0",x"c0",x"a4",x"ac",x"d4",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d0",x"ac",x"8c",x"68",x"64",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"60",x"ac",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"d0",x"ac",x"ac",x"8c",x"6c",x"6c",x"88",x"84",x"80",x"a0",x"a0",x"a0",x"84",x"ac",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"b0",x"b0",x"8c",x"8c",x"88",x"88",x"68",x"48",x"44",x"40",x"60",x"60",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"88",x"ac",x"b0",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"ac",x"ac",x"ac",x"88",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"64",x"88",x"8c",x"ac",x"b0",x"b0",x"b0",x"d0",x"d4",x"f4",x"f9",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f0",x"d0",x"d0",x"d0",x"d0",x"d0",x"d0",x"d0",x"d0",x"d0",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f5",x"f5",x"d5",x"d4",x"b0",x"8c",x"8c",x"8c",x"8c",x"68",x"64",x"60",x"40",x"40",x"40",x"60",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"20",x"20",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"44",x"48",x"48",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"88",x"68",x"44",x"44",x"20",x"20",x"40",x"60",x"60",x"80",x"80",x"80",x"60",x"20",x"24",x"6d",x"91",x"d2",x"f2",x"e9",x"e4",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"84",x"84",x"64",x"84",x"89",x"89",x"85",x"84",x"64",x"80",x"a0",x"c0",x"e0",x"c0",x"c9",x"f6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"d2",x"84",x"40",x"40",x"a0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"80",x"80",x"80",x"80",x"84",x"69",x"69",x"a4",x"e0",x"e0",x"c0",x"c4",x"d4",x"d8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f9",x"f9",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d0",x"b0",x"8c",x"68",x"84",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"40",x"40",x"88",x"cc",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"b0",x"ac",x"ac",x"8c",x"8c",x"6c",x"68",x"84",x"a0",x"a0",x"80",x"80",x"a4",x"ac",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"b0",x"b0",x"8c",x"8c",x"88",x"88",x"68",x"44",x"44",x"40",x"60",x"80",x"80",x"80",x"80",x"80",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"a0",x"a0",x"a0",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"a0",x"80",x"60",x"60",x"80",x"60",x"40",x"40",x"40",x"40",x"40",x"64",x"8c",x"ac",x"b0",x"d0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"ac",x"ac",x"ac",x"88",x"64",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"64",x"88",x"ac",x"ac",x"b0",x"b0",x"b0",x"d0",x"d4",x"f5",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"fd",x"fe",x"fe",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f8",x"f9",x"f9",x"d5",x"d5",x"b0",x"b0",x"8c",x"8c",x"8c",x"6c",x"68",x"64",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"60",x"40",x"60",x"80",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"40",x"40",x"20",x"20",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"44",x"44",x"44",x"64",x"64",x"64",x"60",x"60",x"40",x"20",x"20",x"40",x"80",x"a0",x"80",x"60",x"40",x"20",x"49",x"6d",x"b2",x"d2",x"ed",x"e9",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"a4",x"84",x"84",x"84",x"84",x"85",x"89",x"69",x"44",x"64",x"80",x"c0",x"e0",x"a0",x"a0",x"cd",x"f6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"ad",x"60",x"40",x"60",x"c0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"80",x"80",x"80",x"80",x"64",x"88",x"a4",x"c4",x"e0",x"e0",x"c4",x"cc",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d0",x"b0",x"8c",x"88",x"84",x"80",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"84",x"ac",x"d0",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"ac",x"ac",x"ac",x"8c",x"8c",x"68",x"88",x"a0",x"a0",x"80",x"80",x"a4",x"ac",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"b0",x"b0",x"8c",x"8c",x"88",x"88",x"68",x"48",x"44",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"40",x"40",x"40",x"40",x"40",x"64",x"88",x"ac",x"b0",x"d0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"ac",x"ac",x"ac",x"88",x"64",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"68",x"8c",x"ac",x"ac",x"ac",x"b0",x"b0",x"d4",x"f5",x"f5",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f8",x"f9",x"f9",x"f5",x"d5",x"b0",x"b0",x"8c",x"8c",x"8c",x"6c",x"68",x"64",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"40",x"44",x"49",x"72",x"b2",x"d2",x"ed",x"e9",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"84",x"84",x"84",x"84",x"a8",x"85",x"65",x"45",x"44",x"80",x"c0",x"c0",x"e0",x"a0",x"a9",x"f6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f2",x"85",x"40",x"60",x"a0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"60",x"60",x"80",x"80",x"84",x"68",x"88",x"e0",x"e0",x"e0",x"e8",x"f4",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d0",x"b0",x"ac",x"88",x"84",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"64",x"88",x"d0",x"f4",x"f4",x"f8",x"f4",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"8c",x"88",x"88",x"64",x"80",x"a0",x"a0",x"84",x"ac",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"8c",x"8c",x"88",x"88",x"68",x"68",x"44",x"60",x"60",x"60",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"80",x"60",x"60",x"a0",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"44",x"68",x"ac",x"b0",x"d0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"d0",x"b0",x"ac",x"ac",x"88",x"88",x"64",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"64",x"88",x"8c",x"ac",x"ac",x"b0",x"b0",x"d0",x"d4",x"f5",x"f9",x"f9",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f9",x"f5",x"d4",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"68",x"44",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"60",x"60",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"60",x"40",x"20",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"20",x"20",x"20",x"60",x"80",x"a0",x"80",x"40",x"20",x"24",x"28",x"4d",x"92",x"d6",x"f2",x"e9",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"a0",x"a4",x"a4",x"88",x"a8",x"a9",x"88",x"64",x"64",x"80",x"c0",x"e0",x"c0",x"a0",x"c9",x"d6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"f6",x"c9",x"60",x"20",x"60",x"c0",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"60",x"60",x"84",x"84",x"68",x"84",x"e0",x"e0",x"e8",x"f0",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f9",x"f9",x"f9",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"ac",x"88",x"88",x"64",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"68",x"b0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d0",x"b0",x"ac",x"ac",x"8c",x"8c",x"88",x"88",x"64",x"80",x"80",x"80",x"84",x"ac",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"8c",x"8c",x"88",x"88",x"68",x"68",x"44",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"64",x"8c",x"b0",x"b0",x"d0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"d0",x"b0",x"b0",x"ac",x"ac",x"88",x"64",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"64",x"88",x"8c",x"8c",x"ac",x"b0",x"b0",x"d0",x"d5",x"f9",x"f9",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fd",x"f9",x"f9",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"d4",x"d4",x"d5",x"d4",x"b4",x"b0",x"8c",x"8c",x"8c",x"8c",x"68",x"68",x"44",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"80",x"80",x"60",x"44",x"28",x"4d",x"6d",x"92",x"d2",x"f2",x"ed",x"e5",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a4",x"a4",x"88",x"88",x"88",x"64",x"64",x"80",x"c0",x"c0",x"c0",x"c0",x"c9",x"d2",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"d2",x"84",x"40",x"40",x"80",x"e0",x"e0",x"e0",x"c0",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"84",x"84",x"84",x"a4",x"e0",x"e4",x"ec",x"f4",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fd",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"d4",x"f4",x"f0",x"d0",x"8c",x"88",x"88",x"64",x"60",x"60",x"60",x"60",x"40",x"40",x"64",x"ac",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"b0",x"b0",x"ac",x"8c",x"8c",x"6c",x"68",x"84",x"80",x"80",x"80",x"84",x"a8",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"b0",x"b0",x"8c",x"8c",x"8c",x"88",x"68",x"68",x"64",x"60",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"60",x"60",x"80",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"64",x"88",x"ac",x"b0",x"d0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"d0",x"b0",x"b0",x"ac",x"ac",x"8c",x"64",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"44",x"64",x"88",x"8c",x"8c",x"ac",x"b0",x"b0",x"d4",x"f5",x"f5",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"b4",x"b0",x"90",x"8c",x"8c",x"8c",x"68",x"68",x"44",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"60",x"60",x"a0",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"a0",x"60",x"60",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"40",x"60",x"60",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"60",x"80",x"a0",x"80",x"60",x"40",x"24",x"49",x"71",x"b2",x"d6",x"f6",x"f2",x"e9",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a4",x"84",x"a4",x"a4",x"a4",x"a5",x"89",x"68",x"64",x"64",x"a4",x"c0",x"e0",x"c0",x"a0",x"c9",x"d6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"ad",x"40",x"40",x"80",x"a0",x"e0",x"e0",x"e0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"64",x"68",x"64",x"a4",x"c4",x"e4",x"ec",x"f4",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"fd",x"fd",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f8",x"f8",x"f9",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"f8",x"f8",x"f4",x"f4",x"f4",x"d0",x"b0",x"8c",x"88",x"84",x"64",x"60",x"60",x"60",x"40",x"40",x"60",x"ac",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"b0",x"b0",x"ac",x"ac",x"88",x"6c",x"68",x"84",x"80",x"80",x"80",x"84",x"a8",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"b0",x"b0",x"8c",x"8c",x"8c",x"88",x"68",x"68",x"64",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"88",x"ac",x"b0",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"d4",x"d0",x"b0",x"ac",x"ac",x"ac",x"64",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"44",x"68",x"88",x"8c",x"ac",x"ac",x"b0",x"b0",x"d4",x"d5",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"d4",x"d4",x"b0",x"b0",x"90",x"8c",x"8c",x"8c",x"68",x"68",x"44",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"60",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"80",x"60",x"44",x"49",x"6d",x"92",x"b2",x"d2",x"f2",x"ed",x"e9",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"84",x"84",x"84",x"a4",x"a4",x"a5",x"89",x"69",x"69",x"64",x"a4",x"c0",x"e0",x"e0",x"a0",x"a9",x"d2",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"f2",x"69",x"00",x"40",x"a0",x"c0",x"e0",x"e0",x"e0",x"a0",x"80",x"60",x"80",x"80",x"a0",x"a4",x"85",x"48",x"64",x"c0",x"e0",x"ec",x"f4",x"f9",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"f9",x"f9",x"f9",x"f9",x"f9",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"b4",x"b0",x"d0",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"f9",x"f8",x"f4",x"f4",x"f4",x"d4",x"b0",x"90",x"8c",x"88",x"64",x"60",x"60",x"60",x"40",x"40",x"40",x"ac",x"d0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"b4",x"b0",x"ac",x"8c",x"88",x"88",x"68",x"64",x"64",x"80",x"80",x"84",x"a8",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"8c",x"8c",x"8c",x"8c",x"68",x"68",x"64",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"60",x"60",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"88",x"ac",x"b0",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"d0",x"b0",x"ac",x"b0",x"ac",x"88",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"44",x"68",x"8c",x"8c",x"ac",x"ac",x"b0",x"b0",x"d0",x"d4",x"f5",x"f5",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"b0",x"b0",x"90",x"8c",x"8c",x"8c",x"8c",x"68",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"80",x"a0",x"a0",x"80",x"60",x"40",x"45",x"4d",x"92",x"b6",x"d6",x"f2",x"ee",x"e9",x"e5",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"84",x"64",x"68",x"88",x"a8",x"a9",x"89",x"69",x"49",x"65",x"a4",x"c0",x"e0",x"c0",x"a0",x"a8",x"b2",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"ad",x"64",x"20",x"60",x"c0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"84",x"85",x"65",x"64",x"84",x"e4",x"e8",x"f4",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"f9",x"f9",x"f9",x"f9",x"f5",x"d5",x"d4",x"d4",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"d0",x"d0",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"f9",x"f8",x"f4",x"d4",x"d4",x"b0",x"b0",x"8c",x"88",x"68",x"64",x"64",x"60",x"40",x"40",x"60",x"88",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"b0",x"ac",x"8c",x"8c",x"8c",x"68",x"68",x"64",x"80",x"80",x"80",x"a8",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"b0",x"b0",x"8c",x"8c",x"8c",x"88",x"68",x"64",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"64",x"ac",x"b0",x"d0",x"d0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"b0",x"ac",x"88",x"64",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"64",x"68",x"88",x"8c",x"ac",x"ac",x"8c",x"b0",x"b0",x"d4",x"d5",x"f5",x"f5",x"f5",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"d4",x"d4",x"d0",x"b0",x"b0",x"b0",x"90",x"8c",x"8c",x"6c",x"6c",x"68",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"64",x"69",x"6d",x"72",x"b2",x"d6",x"f2",x"f2",x"ed",x"e9",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"84",x"84",x"88",x"88",x"89",x"89",x"89",x"69",x"69",x"69",x"84",x"c0",x"c0",x"c0",x"c0",x"a8",x"d2",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"d6",x"68",x"40",x"40",x"80",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"84",x"64",x"65",x"65",x"a0",x"c4",x"e8",x"f0",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"f9",x"f9",x"f9",x"f5",x"f5",x"d5",x"b0",x"b0",x"90",x"90",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"ac",x"b0",x"b0",x"b0",x"b0",x"b0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"f9",x"f8",x"d4",x"d4",x"d0",x"d0",x"b0",x"8c",x"68",x"68",x"64",x"44",x"40",x"40",x"60",x"84",x"ac",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"b0",x"ac",x"8c",x"8c",x"8c",x"8c",x"88",x"64",x"60",x"60",x"60",x"84",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"88",x"88",x"64",x"64",x"40",x"60",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"20",x"64",x"88",x"b0",x"d0",x"d0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"d4",x"d4",x"f4",x"f4",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"d0",x"b0",x"b0",x"ac",x"8c",x"88",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"64",x"88",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"d5",x"d5",x"f5",x"f9",x"f9",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"d0",x"d0",x"b0",x"b0",x"8c",x"8c",x"8c",x"6c",x"6c",x"6c",x"68",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"40",x"60",x"80",x"80",x"80",x"a0",x"80",x"40",x"45",x"4d",x"72",x"96",x"da",x"f6",x"f2",x"ed",x"e9",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a4",x"84",x"84",x"84",x"a8",x"a9",x"a9",x"89",x"69",x"48",x"68",x"84",x"a0",x"c0",x"c0",x"a0",x"a9",x"d2",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"d2",x"44",x"40",x"60",x"a0",x"e0",x"e0",x"e0",x"c0",x"80",x"80",x"80",x"80",x"60",x"84",x"84",x"65",x"65",x"a0",x"e4",x"ec",x"f4",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"f9",x"f9",x"f9",x"f5",x"d5",x"d0",x"b0",x"b0",x"8c",x"8c",x"8c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"68",x"68",x"68",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"f9",x"d4",x"d4",x"d4",x"d0",x"b0",x"8c",x"8c",x"68",x"68",x"64",x"40",x"40",x"60",x"84",x"a8",x"d0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"ac",x"8c",x"8c",x"8c",x"8c",x"88",x"64",x"64",x"60",x"60",x"84",x"b0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f9",x"f8",x"f8",x"f4",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"88",x"88",x"88",x"64",x"40",x"60",x"80",x"80",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"20",x"44",x"88",x"ac",x"d0",x"d0",x"d0",x"d0",x"d0",x"d4",x"f4",x"f8",x"f8",x"d4",x"d4",x"f4",x"f4",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"d0",x"b0",x"b0",x"b0",x"8c",x"88",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"68",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"d4",x"d5",x"d5",x"f5",x"f5",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"d0",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"6c",x"6c",x"68",x"48",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"64",x"64",x"69",x"6d",x"6e",x"92",x"b6",x"d6",x"f6",x"f1",x"e9",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a4",x"84",x"84",x"88",x"a9",x"a9",x"89",x"89",x"69",x"68",x"84",x"a4",x"c0",x"c0",x"c0",x"c0",x"c9",x"d2",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"fb",x"b2",x"24",x"40",x"80",x"c0",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"64",x"84",x"84",x"64",x"64",x"c0",x"e8",x"f4",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"fd",x"f9",x"f9",x"f9",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"8c",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"68",x"68",x"68",x"6c",x"6c",x"6c",x"6c",x"8c",x"b0",x"b0",x"b0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"f9",x"f8",x"f4",x"d4",x"d0",x"b0",x"8c",x"8c",x"68",x"68",x"64",x"60",x"40",x"40",x"64",x"88",x"d0",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"ac",x"8c",x"8c",x"8c",x"8c",x"88",x"64",x"64",x"60",x"60",x"84",x"ac",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"8c",x"88",x"88",x"64",x"40",x"60",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"80",x"60",x"40",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"60",x"80",x"60",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"60",x"40",x"40",x"60",x"60",x"40",x"20",x"20",x"40",x"68",x"ac",x"d0",x"d0",x"d0",x"d0",x"d0",x"d4",x"f4",x"f8",x"f8",x"f4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"d0",x"b0",x"b0",x"b0",x"8c",x"88",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"44",x"44",x"68",x"88",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d0",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"68",x"44",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"60",x"60",x"60",x"80",x"60",x"60",x"60",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"40",x"40",x"40",x"60",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"45",x"49",x"4d",x"72",x"b6",x"d6",x"d6",x"f2",x"f2",x"ed",x"e5",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a4",x"84",x"84",x"88",x"a9",x"a9",x"a9",x"a9",x"69",x"69",x"68",x"84",x"c0",x"e0",x"e0",x"c0",x"a0",x"c9",x"f2",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"f6",x"8d",x"24",x"40",x"a0",x"e0",x"e0",x"e0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"64",x"84",x"84",x"60",x"84",x"c4",x"ec",x"f4",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"d5",x"d4",x"b0",x"b0",x"8c",x"8c",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"48",x"68",x"68",x"68",x"68",x"68",x"6c",x"8c",x"8c",x"ac",x"b0",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"f9",x"f8",x"d4",x"d0",x"b0",x"b0",x"8c",x"8c",x"68",x"64",x"64",x"40",x"40",x"60",x"88",x"b0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"8c",x"8c",x"8c",x"8c",x"88",x"64",x"64",x"60",x"60",x"64",x"ac",x"b0",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f4",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"8c",x"88",x"68",x"64",x"44",x"60",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"20",x"40",x"64",x"8c",x"d0",x"d0",x"d0",x"d0",x"d0",x"d4",x"d4",x"f8",x"f8",x"f4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"b0",x"b0",x"b0",x"8c",x"64",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"44",x"68",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"b0",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"b0",x"b0",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"68",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"64",x"64",x"69",x"69",x"8d",x"92",x"96",x"b6",x"d6",x"f2",x"ed",x"ed",x"e9",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a4",x"84",x"84",x"89",x"a9",x"a9",x"a9",x"89",x"69",x"69",x"88",x"a4",x"c0",x"e0",x"e0",x"e0",x"c4",x"cd",x"f6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"db",x"ce",x"65",x"00",x"40",x"c0",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"80",x"64",x"64",x"64",x"80",x"a4",x"ec",x"f4",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f5",x"d4",x"d0",x"b0",x"8c",x"8c",x"6c",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"44",x"44",x"44",x"48",x"44",x"64",x"48",x"48",x"48",x"68",x"68",x"88",x"8c",x"8c",x"b0",x"b0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"f8",x"f4",x"d4",x"b0",x"b0",x"8c",x"8c",x"88",x"68",x"64",x"40",x"40",x"40",x"64",x"ac",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"b0",x"ac",x"8c",x"8c",x"8c",x"88",x"68",x"64",x"60",x"60",x"64",x"88",x"b0",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f4",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"d0",x"b0",x"ac",x"8c",x"8c",x"88",x"68",x"64",x"64",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"60",x"60",x"60",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"60",x"80",x"60",x"40",x"60",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"60",x"60",x"60",x"40",x"40",x"60",x"40",x"20",x"20",x"44",x"88",x"b0",x"b0",x"d0",x"d0",x"d0",x"d0",x"d4",x"f4",x"f8",x"f4",x"f4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"b0",x"b0",x"b0",x"8c",x"64",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"20",x"20",x"40",x"40",x"40",x"44",x"68",x"68",x"8c",x"8c",x"8c",x"8c",x"8c",x"ac",x"b0",x"b0",x"d0",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d0",x"b0",x"b0",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"88",x"68",x"64",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"80",x"a0",x"a0",x"80",x"60",x"60",x"64",x"64",x"69",x"6d",x"8d",x"b2",x"b2",x"d6",x"d7",x"d6",x"ed",x"e9",x"e5",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"84",x"84",x"88",x"89",x"a9",x"a9",x"a9",x"89",x"69",x"49",x"88",x"a4",x"e0",x"e0",x"c0",x"c0",x"c0",x"c9",x"f6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"db",x"a9",x"60",x"00",x"40",x"e0",x"e0",x"e0",x"c0",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"44",x"64",x"a0",x"c4",x"f0",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"f9",x"f9",x"f9",x"f9",x"d5",x"d0",x"b0",x"b0",x"8c",x"8c",x"6c",x"68",x"68",x"48",x"48",x"68",x"68",x"68",x"68",x"68",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"40",x"40",x"40",x"44",x"44",x"44",x"44",x"44",x"64",x"68",x"68",x"88",x"8c",x"ac",x"b0",x"d0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"f8",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"88",x"88",x"64",x"60",x"40",x"40",x"64",x"8c",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"d0",x"ac",x"8c",x"8c",x"8c",x"88",x"68",x"64",x"60",x"60",x"60",x"88",x"ac",x"d0",x"d4",x"d4",x"d4",x"f4",x"f4",x"f8",x"f4",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"88",x"88",x"68",x"64",x"60",x"60",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"88",x"ac",x"b0",x"d0",x"d0",x"d0",x"d0",x"d4",x"f4",x"f8",x"f8",x"f4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"b0",x"b0",x"ac",x"88",x"64",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"20",x"20",x"20",x"40",x"44",x"68",x"68",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"b0",x"d0",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d0",x"b0",x"b0",x"b0",x"b0",x"90",x"8c",x"8c",x"8c",x"8c",x"8c",x"68",x"68",x"68",x"64",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"64",x"64",x"68",x"69",x"8d",x"8d",x"b1",x"b2",x"d2",x"d2",x"ee",x"ee",x"ed",x"e9",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a4",x"a4",x"89",x"89",x"89",x"a9",x"a9",x"a9",x"6d",x"69",x"68",x"84",x"c4",x"c0",x"e0",x"c0",x"c0",x"a9",x"cd",x"d6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"d6",x"85",x"40",x"20",x"60",x"e0",x"e0",x"e0",x"a0",x"80",x"60",x"60",x"60",x"80",x"80",x"80",x"44",x"44",x"c4",x"e8",x"f8",x"fc",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"f9",x"f9",x"f5",x"d4",x"d4",x"b0",x"8c",x"8c",x"8c",x"68",x"68",x"48",x"48",x"48",x"48",x"48",x"68",x"48",x"44",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"44",x"64",x"68",x"88",x"8c",x"ac",x"b0",x"b0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"fd",x"fd",x"f8",x"f8",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"88",x"88",x"64",x"40",x"40",x"40",x"88",x"ac",x"d0",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"d0",x"ac",x"ac",x"8c",x"8c",x"88",x"68",x"64",x"60",x"60",x"60",x"64",x"8c",x"d0",x"d4",x"d0",x"d4",x"f4",x"f4",x"f8",x"f4",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"ac",x"8c",x"8c",x"88",x"68",x"64",x"60",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"60",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"60",x"60",x"40",x"40",x"60",x"80",x"60",x"40",x"60",x"60",x"60",x"60",x"40",x"60",x"60",x"60",x"40",x"60",x"60",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"20",x"20",x"40",x"68",x"ac",x"b0",x"d0",x"d0",x"d0",x"d0",x"d4",x"f4",x"f8",x"f9",x"f4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"d0",x"b0",x"b0",x"b0",x"ac",x"88",x"64",x"60",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"44",x"64",x"68",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"b0",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d0",x"b0",x"b0",x"b0",x"b0",x"90",x"8c",x"8c",x"8c",x"8c",x"6c",x"6c",x"68",x"68",x"68",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"20",x"20",x"20",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"64",x"44",x"49",x"6d",x"6d",x"91",x"b2",x"d2",x"d2",x"f2",x"f2",x"ed",x"e9",x"e5",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a4",x"84",x"84",x"88",x"89",x"a9",x"ad",x"ad",x"8d",x"a9",x"89",x"69",x"68",x"84",x"a4",x"e0",x"e0",x"c0",x"a0",x"a9",x"b2",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"d6",x"44",x"20",x"40",x"80",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"60",x"60",x"60",x"80",x"80",x"40",x"40",x"c8",x"f0",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f5",x"d4",x"d0",x"b0",x"8c",x"8c",x"8c",x"68",x"68",x"48",x"48",x"48",x"48",x"48",x"48",x"44",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"64",x"68",x"68",x"8c",x"8c",x"b0",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"fd",x"fc",x"f8",x"f4",x"d0",x"b0",x"b0",x"ac",x"8c",x"8c",x"88",x"64",x"40",x"20",x"40",x"64",x"ac",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d0",x"d0",x"b0",x"ac",x"8c",x"8c",x"88",x"68",x"64",x"64",x"40",x"40",x"64",x"88",x"d0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"d0",x"ac",x"ac",x"8c",x"8c",x"88",x"68",x"68",x"64",x"60",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"60",x"60",x"60",x"60",x"40",x"60",x"60",x"60",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"60",x"60",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"64",x"88",x"b0",x"d0",x"d0",x"d0",x"d4",x"d4",x"f4",x"f8",x"f9",x"f8",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"b0",x"b0",x"b0",x"ac",x"88",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"40",x"44",x"64",x"68",x"68",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"d0",x"d0",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"b0",x"b0",x"b0",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"6c",x"6c",x"68",x"68",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"64",x"64",x"85",x"89",x"89",x"89",x"8d",x"8d",x"92",x"b2",x"b2",x"d2",x"d2",x"f2",x"ed",x"ed",x"e9",x"e9",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a4",x"a4",x"84",x"89",x"89",x"89",x"ad",x"ad",x"ad",x"8d",x"8d",x"8d",x"89",x"a4",x"c4",x"c0",x"c0",x"a0",x"a0",x"a4",x"cd",x"d6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"fb",x"b2",x"20",x"20",x"60",x"a0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"60",x"60",x"60",x"84",x"80",x"40",x"60",x"cc",x"f4",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f5",x"d4",x"b0",x"b0",x"8c",x"8c",x"88",x"68",x"68",x"68",x"48",x"48",x"48",x"48",x"48",x"44",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"64",x"68",x"88",x"8c",x"b0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fd",x"fc",x"f8",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"88",x"68",x"44",x"40",x"40",x"64",x"88",x"d0",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d0",x"d0",x"ac",x"8c",x"8c",x"88",x"68",x"64",x"64",x"40",x"40",x"40",x"88",x"b0",x"d0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"8c",x"68",x"68",x"64",x"40",x"60",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"60",x"60",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"60",x"60",x"60",x"40",x"40",x"60",x"60",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"44",x"88",x"ac",x"d0",x"b0",x"b0",x"d4",x"d4",x"f4",x"f4",x"f9",x"f8",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"d0",x"b0",x"b0",x"b0",x"ac",x"88",x"64",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"40",x"44",x"64",x"68",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"ac",x"ac",x"b0",x"b0",x"b0",x"b0",x"b0",x"d0",x"d0",x"d0",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d0",x"d0",x"d0",x"d0",x"b0",x"b0",x"b0",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"6c",x"6c",x"68",x"68",x"48",x"44",x"40",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"20",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"64",x"64",x"64",x"69",x"89",x"8d",x"8d",x"92",x"b2",x"b2",x"d6",x"d6",x"f6",x"f2",x"f2",x"ee",x"ed",x"e9",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a4",x"a4",x"84",x"84",x"84",x"89",x"89",x"ad",x"ad",x"ad",x"ad",x"ad",x"8d",x"8d",x"89",x"a8",x"e0",x"e0",x"e0",x"c0",x"a0",x"a4",x"cd",x"d6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"f7",x"ae",x"00",x"20",x"80",x"c0",x"e0",x"e0",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"64",x"60",x"84",x"f0",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f4",x"d4",x"d0",x"b0",x"8c",x"8c",x"8c",x"68",x"68",x"68",x"68",x"48",x"48",x"48",x"44",x"44",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"64",x"68",x"8c",x"ac",x"b0",x"d0",x"d4",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"8c",x"68",x"64",x"40",x"40",x"40",x"88",x"b0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d0",x"d0",x"b0",x"ac",x"8c",x"8c",x"68",x"68",x"64",x"44",x"40",x"40",x"64",x"ac",x"d0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"8c",x"8c",x"68",x"64",x"60",x"40",x"40",x"40",x"60",x"40",x"40",x"60",x"60",x"60",x"60",x"40",x"40",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"60",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"64",x"ac",x"d0",x"b0",x"b0",x"d4",x"d4",x"d4",x"f4",x"f9",x"f8",x"f4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"b0",x"b0",x"ac",x"88",x"64",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"20",x"20",x"20",x"40",x"40",x"44",x"68",x"68",x"88",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"90",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"68",x"68",x"68",x"68",x"44",x"44",x"40",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"64",x"68",x"88",x"89",x"8d",x"8d",x"91",x"b1",x"b2",x"b2",x"b2",x"d2",x"d2",x"d2",x"d2",x"f2",x"ee",x"ed",x"ed",x"e9",x"e5",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a4",x"84",x"84",x"84",x"84",x"a5",x"a9",x"c9",x"cd",x"ad",x"8d",x"8d",x"6d",x"69",x"69",x"88",x"c5",x"e4",x"e0",x"e0",x"c0",x"a0",x"ad",x"d2",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"f2",x"a9",x"00",x"20",x"c0",x"e0",x"e0",x"c0",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"64",x"84",x"a8",x"f4",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f8",x"f4",x"d4",x"d0",x"b0",x"8c",x"8c",x"8c",x"8c",x"68",x"68",x"68",x"48",x"48",x"44",x"44",x"44",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"64",x"68",x"8c",x"ac",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"d0",x"d0",x"ac",x"ac",x"8c",x"8c",x"68",x"68",x"44",x"40",x"40",x"64",x"ac",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d0",x"d0",x"b0",x"ac",x"8c",x"8c",x"68",x"68",x"64",x"44",x"40",x"20",x"64",x"8c",x"b0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"b0",x"ac",x"ac",x"8c",x"8c",x"8c",x"68",x"64",x"60",x"40",x"40",x"40",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"64",x"8c",x"b0",x"b0",x"b0",x"d4",x"d4",x"d4",x"f4",x"f8",x"f8",x"f4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"b0",x"b0",x"b0",x"8c",x"64",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"20",x"20",x"20",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"44",x"44",x"68",x"68",x"68",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"68",x"68",x"68",x"44",x"44",x"44",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"40",x"20",x"20",x"40",x"40",x"40",x"20",x"40",x"40",x"20",x"20",x"40",x"40",x"20",x"20",x"20",x"40",x"40",x"40",x"20",x"20",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"84",x"64",x"64",x"68",x"68",x"69",x"8d",x"91",x"91",x"b2",x"b6",x"d6",x"d6",x"d6",x"f6",x"f2",x"f2",x"ee",x"ed",x"ed",x"e9",x"e9",x"e5",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"e4",x"c4",x"a4",x"84",x"84",x"84",x"89",x"a9",x"a9",x"c9",x"cd",x"ce",x"ad",x"8d",x"8d",x"69",x"89",x"84",x"a4",x"e0",x"e0",x"e0",x"c0",x"a0",x"a9",x"d6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"fb",x"ee",x"85",x"00",x"20",x"c0",x"e0",x"e0",x"c0",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"64",x"88",x"d0",x"f4",x"f8",x"fc",x"fc",x"f8",x"f8",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"8c",x"6c",x"68",x"68",x"68",x"48",x"44",x"44",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"64",x"68",x"8c",x"ac",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d0",x"d0",x"ac",x"ac",x"8c",x"8c",x"68",x"68",x"44",x"40",x"40",x"64",x"ac",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f0",x"d0",x"b0",x"ac",x"8c",x"8c",x"68",x"68",x"68",x"44",x"40",x"20",x"44",x"88",x"b0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"d0",x"b0",x"ac",x"8c",x"8c",x"8c",x"8c",x"68",x"64",x"60",x"60",x"40",x"40",x"40",x"60",x"60",x"60",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"60",x"60",x"60",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"44",x"8c",x"b0",x"b0",x"b0",x"d4",x"d4",x"d4",x"f4",x"f4",x"f8",x"f4",x"f4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"b0",x"b0",x"ac",x"64",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"44",x"44",x"68",x"68",x"88",x"8c",x"6c",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"90",x"90",x"90",x"90",x"90",x"90",x"90",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"6c",x"6c",x"6c",x"68",x"68",x"68",x"68",x"68",x"44",x"44",x"44",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"20",x"20",x"40",x"40",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"20",x"20",x"20",x"40",x"20",x"20",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"64",x"64",x"68",x"69",x"6d",x"8d",x"91",x"91",x"b6",x"b6",x"b6",x"d6",x"d6",x"d6",x"d2",x"f2",x"ee",x"ed",x"e9",x"e9",x"e5",x"e5",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a4",x"a4",x"84",x"84",x"a4",x"a5",x"a5",x"a9",x"a9",x"ad",x"ae",x"b2",x"91",x"8d",x"6d",x"89",x"89",x"c5",x"c4",x"e0",x"e0",x"c0",x"c0",x"c0",x"c9",x"d2",x"d6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"fb",x"c9",x"64",x"00",x"40",x"e0",x"e0",x"e0",x"a0",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"40",x"44",x"8c",x"d4",x"f8",x"f8",x"fc",x"fd",x"f8",x"f8",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"b0",x"b0",x"8c",x"8c",x"88",x"68",x"68",x"68",x"68",x"68",x"48",x"44",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"20",x"20",x"40",x"40",x"20",x"20",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"64",x"68",x"8c",x"ac",x"b0",x"d0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d0",x"d0",x"b0",x"ac",x"8c",x"68",x"68",x"68",x"64",x"44",x"40",x"40",x"ac",x"d0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f0",x"d0",x"d0",x"ac",x"8c",x"8c",x"6c",x"68",x"68",x"44",x"40",x"20",x"40",x"88",x"ac",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"8c",x"8c",x"68",x"64",x"60",x"60",x"40",x"20",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"40",x"88",x"b0",x"b0",x"b0",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"b0",x"b0",x"ac",x"68",x"64",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"44",x"44",x"68",x"68",x"68",x"68",x"68",x"6c",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"6c",x"6c",x"68",x"68",x"68",x"68",x"68",x"44",x"44",x"44",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"20",x"20",x"40",x"40",x"20",x"20",x"40",x"40",x"40",x"40",x"20",x"40",x"40",x"20",x"20",x"40",x"40",x"20",x"20",x"20",x"40",x"20",x"20",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"84",x"69",x"69",x"6d",x"6d",x"71",x"91",x"96",x"b6",x"d6",x"f6",x"f6",x"f6",x"f2",x"f2",x"f2",x"ed",x"e9",x"e9",x"e5",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c4",x"c4",x"a4",x"a4",x"84",x"89",x"89",x"89",x"a9",x"a9",x"a9",x"ad",x"ad",x"ae",x"b2",x"92",x"8d",x"6d",x"89",x"a4",x"c4",x"e0",x"e0",x"e0",x"e0",x"c0",x"a4",x"a9",x"d2",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"fb",x"a9",x"40",x"00",x"40",x"e0",x"e0",x"e0",x"a0",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"40",x"44",x"8c",x"d4",x"f8",x"f8",x"f9",x"f9",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"68",x"68",x"68",x"68",x"68",x"68",x"44",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"64",x"88",x"ac",x"b0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d0",x"d0",x"ac",x"8c",x"68",x"68",x"68",x"68",x"44",x"20",x"40",x"ac",x"d0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f0",x"d0",x"d0",x"ac",x"8c",x"8c",x"8c",x"68",x"68",x"44",x"40",x"20",x"40",x"68",x"ac",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"8c",x"8c",x"88",x"64",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"68",x"b0",x"b0",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f9",x"f8",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f4",x"d4",x"d0",x"b0",x"b0",x"b0",x"b0",x"ac",x"88",x"64",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"44",x"48",x"48",x"68",x"68",x"68",x"6c",x"6c",x"6c",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"68",x"68",x"44",x"44",x"44",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"80",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"64",x"68",x"68",x"69",x"8d",x"92",x"b2",x"b2",x"b2",x"b6",x"d6",x"d6",x"d6",x"d2",x"f2",x"ee",x"ed",x"e9",x"e9",x"e9",x"e5",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a4",x"a4",x"a4",x"84",x"84",x"a9",x"a9",x"a9",x"a9",x"a9",x"ad",x"cd",x"cd",x"ad",x"92",x"92",x"72",x"6d",x"8d",x"a9",x"c5",x"e1",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a9",x"d2",x"da",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"db",x"85",x"40",x"20",x"60",x"e0",x"e0",x"c0",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"40",x"44",x"b0",x"f8",x"f8",x"f8",x"f9",x"f9",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"68",x"68",x"68",x"68",x"48",x"48",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"64",x"8c",x"ac",x"d0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d0",x"d0",x"ac",x"8c",x"68",x"68",x"68",x"68",x"44",x"20",x"40",x"8c",x"b0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"d0",x"ac",x"8c",x"8c",x"8c",x"68",x"68",x"64",x"40",x"20",x"40",x"64",x"8c",x"d0",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"ac",x"8c",x"8c",x"8c",x"88",x"64",x"44",x"40",x"40",x"60",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"68",x"8c",x"b0",x"d0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f9",x"f8",x"d4",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f4",x"d4",x"d4",x"b0",x"b0",x"b0",x"b0",x"ac",x"88",x"64",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"44",x"44",x"44",x"44",x"44",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"6c",x"68",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"44",x"44",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"20",x"20",x"40",x"40",x"20",x"20",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"40",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"64",x"64",x"68",x"69",x"6d",x"8d",x"91",x"91",x"92",x"b6",x"d6",x"d6",x"d6",x"f6",x"f2",x"f2",x"f2",x"ed",x"ed",x"e9",x"e5",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a4",x"a4",x"a4",x"a4",x"84",x"88",x"88",x"89",x"a9",x"ad",x"ad",x"cd",x"cd",x"cd",x"b2",x"b2",x"92",x"91",x"91",x"8d",x"8d",x"a9",x"c5",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a4",x"a9",x"d6",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"d6",x"44",x"40",x"60",x"a0",x"e0",x"e0",x"a0",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"64",x"88",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"8c",x"88",x"68",x"68",x"48",x"48",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"68",x"8c",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d0",x"d0",x"ac",x"8c",x"88",x"68",x"68",x"68",x"44",x"40",x"40",x"64",x"8c",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"88",x"68",x"68",x"44",x"20",x"20",x"40",x"88",x"b0",x"d0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"8c",x"88",x"68",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"64",x"88",x"b0",x"b0",x"b0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f9",x"f8",x"f4",x"d4",x"d4",x"d4",x"f4",x"f8",x"f8",x"f4",x"d4",x"d4",x"d4",x"b0",x"b0",x"b0",x"b0",x"ac",x"88",x"60",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"44",x"44",x"64",x"68",x"68",x"68",x"68",x"68",x"68",x"6c",x"8c",x"6c",x"6c",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"44",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"44",x"45",x"49",x"69",x"6d",x"91",x"92",x"b2",x"b6",x"d6",x"d6",x"d6",x"d6",x"d6",x"f2",x"f1",x"ed",x"ed",x"e9",x"e9",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c4",x"a4",x"a4",x"84",x"84",x"84",x"84",x"84",x"88",x"89",x"a9",x"a9",x"a9",x"a9",x"cd",x"cd",x"cd",x"cd",x"b2",x"b2",x"91",x"71",x"6d",x"6d",x"8d",x"a9",x"c9",x"e4",x"e4",x"e0",x"c0",x"a0",x"a0",x"a0",x"a4",x"cd",x"d6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"d6",x"44",x"20",x"80",x"c0",x"e0",x"c0",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"84",x"ac",x"f4",x"f8",x"f8",x"f8",x"f8",x"fc",x"f8",x"f8",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"88",x"68",x"68",x"48",x"44",x"24",x"20",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"64",x"88",x"ac",x"b0",x"d0",x"d0",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d0",x"d0",x"ac",x"8c",x"8c",x"88",x"68",x"68",x"44",x"44",x"40",x"40",x"68",x"d0",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"d0",x"ac",x"8c",x"8c",x"88",x"68",x"68",x"44",x"20",x"20",x"20",x"68",x"b0",x"d0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"68",x"64",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"44",x"68",x"ac",x"d0",x"b0",x"b0",x"d4",x"d4",x"f4",x"f8",x"f9",x"f8",x"f4",x"d4",x"d4",x"d4",x"d4",x"f8",x"f8",x"f4",x"d4",x"d4",x"d4",x"d0",x"b0",x"b0",x"b0",x"ac",x"88",x"60",x"40",x"40",x"40",x"60",x"60",x"60",x"40",x"40",x"20",x"20",x"20",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"44",x"44",x"44",x"44",x"44",x"68",x"68",x"68",x"68",x"68",x"68",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"44",x"20",x"20",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"84",x"84",x"84",x"84",x"69",x"4d",x"6d",x"6d",x"92",x"92",x"b6",x"d6",x"d6",x"f6",x"f6",x"f2",x"f2",x"f2",x"ed",x"ed",x"e9",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c4",x"c4",x"c4",x"a5",x"a9",x"89",x"89",x"89",x"89",x"89",x"89",x"89",x"ad",x"ad",x"ad",x"cd",x"ce",x"ce",x"d2",x"b2",x"b2",x"b1",x"b1",x"8d",x"8d",x"89",x"89",x"a5",x"c4",x"e4",x"e0",x"e0",x"c0",x"c0",x"a0",x"a4",x"a9",x"b1",x"d6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"b6",x"24",x"20",x"80",x"c0",x"e0",x"c0",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"84",x"ac",x"f4",x"f8",x"f8",x"f8",x"f8",x"fc",x"f8",x"f8",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"b0",x"ac",x"8c",x"8c",x"8c",x"88",x"68",x"68",x"68",x"48",x"48",x"24",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"20",x"20",x"40",x"40",x"20",x"40",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"20",x"20",x"40",x"60",x"88",x"8c",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d0",x"d0",x"ac",x"8c",x"8c",x"88",x"68",x"68",x"44",x"44",x"40",x"40",x"68",x"b0",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"d0",x"ac",x"ac",x"8c",x"88",x"68",x"68",x"48",x"24",x"20",x"20",x"68",x"ac",x"b0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"b0",x"b0",x"ac",x"8c",x"8c",x"8c",x"68",x"64",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"64",x"ac",x"d0",x"b0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"d4",x"d4",x"d0",x"b0",x"b0",x"b0",x"ac",x"88",x"60",x"40",x"40",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"44",x"44",x"48",x"49",x"6d",x"6d",x"92",x"b2",x"b2",x"d6",x"d6",x"d6",x"d6",x"d2",x"d2",x"f2",x"ed",x"ed",x"e9",x"e9",x"e5",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a4",x"a4",x"a4",x"84",x"84",x"84",x"89",x"a9",x"a9",x"a9",x"a9",x"c9",x"cd",x"ad",x"ad",x"ae",x"ae",x"ce",x"ce",x"d2",x"b2",x"b2",x"92",x"92",x"92",x"91",x"8d",x"8d",x"a9",x"e5",x"e1",x"e1",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a4",x"cd",x"d6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"b2",x"24",x"20",x"80",x"c0",x"e0",x"c0",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"88",x"cc",x"f4",x"f8",x"f8",x"f8",x"f8",x"fc",x"f8",x"f8",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"b0",x"ac",x"8c",x"8c",x"8c",x"88",x"68",x"68",x"68",x"48",x"44",x"24",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"64",x"88",x"ac",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d0",x"d0",x"b0",x"8c",x"8c",x"88",x"68",x"68",x"44",x"44",x"40",x"40",x"64",x"ac",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"d0",x"b0",x"ac",x"8c",x"8c",x"88",x"68",x"68",x"44",x"20",x"20",x"64",x"8c",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"8c",x"88",x"64",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"44",x"8c",x"d0",x"d0",x"d4",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"d4",x"d4",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f4",x"d4",x"d0",x"b0",x"b0",x"b0",x"b0",x"88",x"60",x"40",x"40",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"84",x"84",x"84",x"84",x"64",x"69",x"69",x"6d",x"6d",x"6d",x"91",x"b2",x"b2",x"d6",x"d6",x"f2",x"f2",x"f2",x"f2",x"ed",x"ed",x"e9",x"e9",x"e5",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c4",x"c4",x"a5",x"a5",x"85",x"85",x"89",x"89",x"89",x"89",x"89",x"8d",x"ad",x"ad",x"ad",x"cd",x"cd",x"ce",x"ae",x"ae",x"b2",x"b2",x"b2",x"b2",x"b2",x"b2",x"b2",x"ad",x"ad",x"a9",x"a9",x"a9",x"c5",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c4",x"a4",x"a9",x"d1",x"f6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"fb",x"b2",x"20",x"20",x"a0",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"a8",x"d0",x"f4",x"f8",x"f8",x"f8",x"f8",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"88",x"68",x"68",x"68",x"48",x"48",x"44",x"44",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"20",x"20",x"40",x"64",x"ac",x"b0",x"d0",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"8c",x"8c",x"88",x"68",x"68",x"44",x"44",x"40",x"20",x"44",x"8c",x"b0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"d0",x"b0",x"ac",x"8c",x"8c",x"88",x"68",x"68",x"44",x"20",x"20",x"44",x"88",x"ac",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"ac",x"8c",x"8c",x"88",x"68",x"44",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"8c",x"b0",x"d0",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f4",x"d4",x"d4",x"d4",x"f4",x"f8",x"f9",x"f9",x"f8",x"d4",x"d4",x"b0",x"b0",x"b0",x"b0",x"ac",x"60",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"44",x"44",x"48",x"6d",x"6d",x"8e",x"92",x"b2",x"b2",x"d2",x"d2",x"f2",x"f2",x"f2",x"ed",x"ed",x"ed",x"ed",x"e9",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a4",x"a4",x"84",x"84",x"84",x"89",x"89",x"89",x"a9",x"a9",x"a9",x"a9",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"b1",x"b2",x"b2",x"b2",x"b2",x"b2",x"b2",x"92",x"92",x"92",x"91",x"8d",x"ad",x"c9",x"c5",x"e5",x"e1",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"a0",x"a9",x"f2",x"f6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"fa",x"b2",x"20",x"20",x"a0",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"64",x"ac",x"d0",x"f4",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"8c",x"8c",x"8c",x"68",x"68",x"68",x"68",x"48",x"48",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"40",x"20",x"20",x"40",x"64",x"8c",x"b0",x"d0",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"8c",x"8c",x"88",x"68",x"68",x"44",x"44",x"40",x"20",x"44",x"8c",x"b0",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"8c",x"88",x"68",x"44",x"40",x"20",x"44",x"68",x"8c",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"ac",x"8c",x"8c",x"8c",x"68",x"64",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"88",x"b0",x"d0",x"d4",x"d0",x"d4",x"d4",x"f4",x"f4",x"f9",x"f9",x"f4",x"d4",x"d4",x"d4",x"f4",x"f9",x"f9",x"f9",x"f4",x"d4",x"d4",x"b0",x"b0",x"b0",x"b0",x"ac",x"60",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"84",x"84",x"84",x"84",x"85",x"69",x"69",x"6d",x"6d",x"6d",x"92",x"92",x"b2",x"b2",x"d2",x"f2",x"f2",x"ee",x"ee",x"ed",x"e9",x"e9",x"e9",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a4",x"a4",x"a4",x"a4",x"84",x"84",x"89",x"89",x"89",x"89",x"89",x"8d",x"8d",x"ad",x"ad",x"ad",x"ad",x"ad",x"ae",x"b2",x"b2",x"b2",x"b2",x"b2",x"b2",x"b2",x"b2",x"b2",x"b2",x"ad",x"ad",x"ad",x"ad",x"ad",x"a9",x"a9",x"c5",x"c4",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a4",x"a4",x"a9",x"ad",x"d2",x"fa",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"f6",x"8d",x"00",x"20",x"a0",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"84",x"ac",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"8c",x"8c",x"88",x"68",x"68",x"68",x"68",x"48",x"44",x"24",x"44",x"40",x"40",x"40",x"40",x"60",x"40",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"20",x"20",x"40",x"20",x"44",x"88",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"88",x"68",x"68",x"68",x"44",x"40",x"20",x"40",x"68",x"ac",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"d0",x"b0",x"ac",x"8c",x"8c",x"88",x"68",x"68",x"44",x"20",x"40",x"64",x"8c",x"b0",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"ac",x"ac",x"8c",x"8c",x"88",x"88",x"40",x"20",x"60",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"68",x"ac",x"b0",x"d4",x"b0",x"d4",x"d4",x"f4",x"f4",x"f9",x"f9",x"f8",x"d4",x"d4",x"d4",x"d4",x"f8",x"f9",x"f9",x"f4",x"d4",x"d4",x"b0",x"b0",x"b0",x"b0",x"ac",x"60",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"60",x"40",x"64",x"64",x"69",x"6d",x"6d",x"71",x"91",x"92",x"b2",x"b2",x"d2",x"d2",x"d2",x"d2",x"ce",x"ee",x"ed",x"e9",x"e9",x"e5",x"e5",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a4",x"a4",x"84",x"84",x"84",x"84",x"84",x"84",x"88",x"89",x"89",x"89",x"89",x"ad",x"ad",x"ad",x"ce",x"ce",x"ce",x"cd",x"ad",x"b1",x"b1",x"b2",x"b2",x"b2",x"92",x"92",x"92",x"92",x"b2",x"b2",x"b2",x"b2",x"ad",x"cd",x"c9",x"e9",x"e5",x"e4",x"e0",x"e0",x"e0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"88",x"91",x"d6",x"da",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"f2",x"8d",x"00",x"20",x"c0",x"e0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"84",x"cc",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"8c",x"8c",x"68",x"68",x"68",x"68",x"68",x"48",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"20",x"40",x"68",x"ac",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"88",x"68",x"68",x"68",x"44",x"44",x"20",x"20",x"68",x"8c",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"d0",x"b0",x"ac",x"8c",x"8c",x"8c",x"68",x"68",x"44",x"20",x"20",x"44",x"88",x"b0",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"ac",x"8c",x"8c",x"8c",x"88",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"64",x"8c",x"b0",x"d4",x"d0",x"d4",x"d4",x"d4",x"f4",x"f9",x"f9",x"f9",x"f4",x"d4",x"d4",x"d4",x"f4",x"f9",x"f5",x"d4",x"d4",x"d0",x"b0",x"b0",x"b0",x"b0",x"8c",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"84",x"84",x"84",x"84",x"85",x"89",x"89",x"8d",x"8d",x"91",x"92",x"b2",x"b2",x"d2",x"d2",x"ce",x"ee",x"ee",x"ed",x"e9",x"e9",x"e9",x"e5",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a4",x"a4",x"a4",x"84",x"84",x"84",x"84",x"89",x"89",x"89",x"a9",x"a9",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ae",x"ae",x"ae",x"b2",x"b2",x"91",x"b1",x"b1",x"b1",x"b1",x"b1",x"b1",x"ad",x"ad",x"ad",x"a9",x"c9",x"c9",x"c9",x"c9",x"c4",x"c4",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"84",x"a8",x"a8",x"a9",x"ad",x"b6",x"da",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"d2",x"8d",x"00",x"20",x"c0",x"e0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"d0",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"8c",x"8c",x"68",x"68",x"68",x"68",x"48",x"48",x"44",x"44",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"60",x"60",x"60",x"40",x"60",x"60",x"60",x"60",x"40",x"40",x"60",x"40",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"40",x"68",x"8c",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"88",x"68",x"68",x"68",x"44",x"44",x"20",x"20",x"44",x"88",x"b0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"8c",x"88",x"68",x"44",x"20",x"20",x"20",x"68",x"b0",x"d0",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"ac",x"ac",x"8c",x"8c",x"68",x"64",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"44",x"68",x"b0",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"f9",x"f9",x"f9",x"f4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"b0",x"b0",x"b0",x"b0",x"ac",x"88",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"60",x"60",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"40",x"44",x"44",x"49",x"49",x"49",x"4d",x"6d",x"b2",x"b2",x"b2",x"d2",x"d2",x"d2",x"ee",x"ed",x"ed",x"e9",x"e9",x"e5",x"e5",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a9",x"89",x"89",x"a9",x"ad",x"ad",x"cd",x"cd",x"cd",x"cd",x"ce",x"ce",x"b2",x"b2",x"b1",x"91",x"91",x"91",x"71",x"71",x"92",x"91",x"91",x"91",x"ad",x"ad",x"cd",x"c9",x"c9",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"60",x"60",x"60",x"64",x"89",x"ad",x"d2",x"fa",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"d2",x"89",x"00",x"20",x"c0",x"e0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"88",x"d0",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"8c",x"8c",x"68",x"68",x"68",x"68",x"44",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"40",x"64",x"8c",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"88",x"68",x"68",x"68",x"48",x"44",x"20",x"20",x"44",x"68",x"ac",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"ac",x"8c",x"8c",x"8c",x"68",x"68",x"44",x"20",x"20",x"68",x"ac",x"b0",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"ac",x"ac",x"8c",x"8c",x"88",x"64",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"44",x"b0",x"d5",x"d4",x"d4",x"d4",x"d4",x"d4",x"f5",x"f9",x"f9",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"b0",x"b0",x"b0",x"b0",x"b0",x"8c",x"8c",x"68",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"64",x"64",x"64",x"64",x"64",x"68",x"69",x"69",x"6d",x"6d",x"8d",x"6d",x"6d",x"ae",x"d2",x"cd",x"cd",x"cd",x"e9",x"e9",x"e9",x"e5",x"e5",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a4",x"a5",x"a9",x"a9",x"a9",x"a9",x"a9",x"ad",x"ad",x"ad",x"ae",x"ae",x"ae",x"ad",x"ad",x"b2",x"b2",x"b1",x"b1",x"b1",x"b1",x"b1",x"ad",x"8d",x"8d",x"ad",x"ad",x"ad",x"a9",x"c9",x"c9",x"c5",x"c4",x"c4",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"84",x"84",x"88",x"89",x"8d",x"b1",x"b6",x"d6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ce",x"89",x"00",x"20",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"88",x"d0",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"8c",x"8c",x"68",x"68",x"68",x"68",x"44",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"60",x"80",x"40",x"40",x"60",x"80",x"60",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"60",x"40",x"20",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"44",x"88",x"b0",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"b0",x"ac",x"8c",x"88",x"68",x"68",x"68",x"68",x"44",x"20",x"20",x"40",x"68",x"ac",x"b0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"8c",x"6c",x"68",x"44",x"20",x"20",x"64",x"8c",x"b0",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"ac",x"8c",x"68",x"44",x"60",x"40",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"44",x"8c",x"d1",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"f5",x"d5",x"d4",x"d4",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"8c",x"8c",x"68",x"64",x"40",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"40",x"40",x"44",x"48",x"48",x"49",x"69",x"6d",x"8d",x"ad",x"ad",x"cd",x"cd",x"cd",x"cd",x"cd",x"cd",x"ed",x"e9",x"e9",x"e5",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a4",x"a4",x"84",x"84",x"84",x"85",x"a5",x"a5",x"a9",x"a9",x"a9",x"a9",x"a9",x"a9",x"ad",x"ad",x"ad",x"ae",x"b2",x"b2",x"b2",x"ae",x"ad",x"8d",x"91",x"91",x"91",x"91",x"91",x"91",x"ad",x"ad",x"cd",x"c9",x"c9",x"c9",x"e5",x"e5",x"e5",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"60",x"60",x"60",x"84",x"88",x"89",x"ad",x"b2",x"d6",x"da",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ce",x"89",x"00",x"20",x"c0",x"c0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"88",x"d0",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"8c",x"8c",x"68",x"68",x"68",x"68",x"44",x"44",x"24",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"44",x"68",x"b0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"b0",x"ac",x"8c",x"88",x"68",x"68",x"68",x"68",x"44",x"20",x"20",x"20",x"44",x"8c",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"8c",x"6c",x"68",x"44",x"20",x"20",x"44",x"8c",x"b0",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"90",x"8c",x"8c",x"8c",x"88",x"64",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"68",x"b0",x"b0",x"d4",x"b0",x"b0",x"b0",x"d4",x"d4",x"d4",x"d4",x"b0",x"b0",x"b0",x"b0",x"b0",x"90",x"90",x"90",x"90",x"8c",x"8c",x"68",x"64",x"44",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"64",x"64",x"64",x"68",x"68",x"69",x"69",x"69",x"8d",x"8d",x"8d",x"ad",x"ad",x"cd",x"cd",x"ed",x"ed",x"e9",x"e9",x"e9",x"e9",x"e5",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a4",x"a4",x"84",x"84",x"84",x"84",x"88",x"88",x"89",x"a9",x"a9",x"a9",x"a9",x"a9",x"ad",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"91",x"92",x"b2",x"b1",x"8d",x"8d",x"8d",x"ad",x"ad",x"ad",x"ad",x"c9",x"c9",x"c9",x"c5",x"c4",x"c4",x"e4",x"e0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a4",x"a4",x"a5",x"a9",x"a9",x"ad",x"ad",x"b2",x"b2",x"d6",x"d6",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"cd",x"89",x"00",x"20",x"c0",x"c0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"84",x"88",x"d0",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"8c",x"8c",x"68",x"68",x"68",x"68",x"44",x"44",x"24",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"60",x"60",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"20",x"40",x"40",x"20",x"20",x"40",x"68",x"b0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"b0",x"ac",x"8c",x"8c",x"68",x"68",x"68",x"68",x"44",x"20",x"20",x"20",x"44",x"88",x"b0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"8c",x"8c",x"8c",x"6c",x"68",x"68",x"40",x"20",x"44",x"68",x"b0",x"b4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"b0",x"b0",x"b0",x"90",x"8c",x"8c",x"88",x"88",x"40",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"20",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"64",x"8c",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"90",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"68",x"68",x"44",x"20",x"20",x"20",x"20",x"20",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"40",x"44",x"24",x"24",x"48",x"48",x"4d",x"6d",x"8d",x"91",x"91",x"cd",x"ed",x"ed",x"ed",x"e9",x"e9",x"e9",x"e9",x"e5",x"e5",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"a4",x"a5",x"84",x"84",x"84",x"84",x"84",x"84",x"88",x"88",x"89",x"89",x"89",x"89",x"89",x"ad",x"ad",x"ad",x"ad",x"ad",x"8d",x"8d",x"91",x"91",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"ad",x"ad",x"c9",x"c9",x"e9",x"e5",x"e4",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"60",x"60",x"64",x"89",x"8d",x"ae",x"d2",x"d6",x"fb",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"cd",x"89",x"00",x"20",x"c0",x"c0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"84",x"a8",x"d0",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"8c",x"8c",x"68",x"68",x"68",x"68",x"44",x"24",x"24",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"40",x"60",x"60",x"60",x"40",x"60",x"60",x"60",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"64",x"b0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"b0",x"ac",x"8c",x"8c",x"68",x"68",x"68",x"68",x"44",x"20",x"20",x"00",x"40",x"88",x"ac",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"d0",x"b0",x"ac",x"8c",x"8c",x"6c",x"68",x"68",x"44",x"20",x"44",x"68",x"90",x"d4",x"d4",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f4",x"f4",x"d4",x"b0",x"b0",x"b0",x"90",x"8c",x"8c",x"8c",x"88",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"68",x"8c",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"90",x"90",x"90",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"68",x"44",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"44",x"44",x"44",x"64",x"69",x"69",x"69",x"89",x"8d",x"ad",x"ad",x"ad",x"cd",x"c9",x"c9",x"e9",x"e9",x"e5",x"e5",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a4",x"a4",x"84",x"84",x"84",x"84",x"84",x"89",x"89",x"89",x"a9",x"a9",x"a9",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"ad",x"ad",x"a9",x"c9",x"c9",x"c9",x"c5",x"c4",x"c4",x"c4",x"c4",x"c4",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a4",x"a9",x"a9",x"a9",x"ad",x"ad",x"b1",x"b2",x"b6",x"d6",x"db",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ad",x"89",x"00",x"20",x"c0",x"c0",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"60",x"84",x"a8",x"d0",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"8c",x"8c",x"68",x"68",x"68",x"68",x"44",x"24",x"24",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"60",x"60",x"60",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"64",x"ac",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"b0",x"ac",x"8c",x"8c",x"68",x"68",x"68",x"68",x"44",x"24",x"20",x"00",x"20",x"68",x"ac",x"b0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"6c",x"68",x"68",x"44",x"20",x"40",x"64",x"8c",x"d4",x"d0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"b0",x"90",x"90",x"8c",x"8c",x"8c",x"88",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"44",x"68",x"8c",x"b0",x"b0",x"b0",x"90",x"90",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"8c",x"8c",x"6c",x"68",x"68",x"44",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"60",x"80",x"a0",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"44",x"24",x"24",x"24",x"24",x"49",x"49",x"69",x"69",x"89",x"ad",x"cd",x"ed",x"e9",x"e9",x"e9",x"e5",x"e5",x"e5",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a4",x"a4",x"84",x"84",x"84",x"84",x"84",x"85",x"85",x"85",x"84",x"84",x"88",x"88",x"a9",x"a9",x"a9",x"a9",x"a9",x"ad",x"ad",x"ad",x"ad",x"ad",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"ad",x"a9",x"c9",x"c9",x"e5",x"e5",x"e1",x"e1",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a0",x"80",x"60",x"60",x"60",x"64",x"84",x"88",x"89",x"ad",x"d2",x"d6",x"d6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ad",x"89",x"00",x"20",x"a0",x"c0",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"84",x"a8",x"d0",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"8c",x"8c",x"68",x"68",x"68",x"68",x"44",x"24",x"24",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"64",x"ac",x"d4",x"d4",x"f4",x"f8",x"f8",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"b0",x"ac",x"8c",x"8c",x"68",x"68",x"68",x"68",x"44",x"44",x"20",x"00",x"20",x"44",x"8c",x"b0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"68",x"44",x"20",x"20",x"44",x"8c",x"b0",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f9",x"f9",x"f8",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f4",x"d4",x"d0",x"b0",x"b0",x"8c",x"ac",x"ac",x"8c",x"8c",x"64",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"44",x"68",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"68",x"68",x"68",x"68",x"48",x"44",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"44",x"44",x"44",x"44",x"48",x"68",x"69",x"69",x"89",x"89",x"89",x"a9",x"a9",x"a9",x"c9",x"c9",x"e9",x"e5",x"e5",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a4",x"a4",x"a4",x"84",x"84",x"84",x"84",x"85",x"89",x"89",x"a9",x"a9",x"89",x"89",x"89",x"89",x"89",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"a9",x"c9",x"c9",x"c9",x"c9",x"c9",x"c4",x"c4",x"c4",x"c4",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"84",x"84",x"84",x"89",x"a9",x"ad",x"ad",x"b2",x"b2",x"d6",x"d6",x"db",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"cd",x"89",x"04",x"20",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"88",x"d0",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"b0",x"ac",x"8c",x"88",x"68",x"68",x"68",x"44",x"24",x"24",x"44",x"40",x"40",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"40",x"68",x"b0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f5",x"d4",x"b0",x"8c",x"8c",x"8c",x"6c",x"68",x"68",x"48",x"44",x"40",x"20",x"20",x"20",x"40",x"68",x"b0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"8c",x"8c",x"68",x"40",x"20",x"20",x"68",x"b0",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f9",x"f9",x"f9",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f4",x"d4",x"d4",x"d0",x"b0",x"ac",x"b0",x"b0",x"90",x"8c",x"68",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"20",x"20",x"20",x"20",x"00",x"00",x"20",x"20",x"44",x"48",x"68",x"6c",x"6c",x"6c",x"8c",x"8c",x"8c",x"8c",x"6c",x"6c",x"68",x"68",x"48",x"48",x"44",x"44",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"44",x"24",x"24",x"24",x"24",x"28",x"28",x"48",x"69",x"69",x"8d",x"ad",x"cd",x"ed",x"e9",x"e9",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"a5",x"a9",x"a9",x"a9",x"a9",x"a9",x"a9",x"a9",x"a9",x"a9",x"ad",x"8d",x"8d",x"8d",x"6d",x"6d",x"6d",x"6d",x"89",x"89",x"89",x"89",x"a9",x"c9",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"40",x"44",x"64",x"69",x"89",x"8d",x"b2",x"d6",x"d6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"cd",x"89",x"04",x"20",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"88",x"d0",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d0",x"d0",x"ac",x"8c",x"88",x"68",x"68",x"68",x"44",x"44",x"24",x"44",x"40",x"40",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"40",x"68",x"b0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f5",x"d4",x"b0",x"8c",x"8c",x"8c",x"6c",x"68",x"68",x"48",x"44",x"40",x"20",x"20",x"20",x"20",x"68",x"b0",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"8c",x"8c",x"68",x"44",x"20",x"20",x"68",x"b0",x"b0",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f9",x"f9",x"f9",x"f8",x"f4",x"f4",x"f4",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"b0",x"b0",x"90",x"8c",x"68",x"64",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"20",x"20",x"20",x"24",x"44",x"48",x"48",x"68",x"68",x"68",x"6c",x"6c",x"6c",x"68",x"68",x"48",x"44",x"24",x"24",x"20",x"20",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"44",x"44",x"44",x"44",x"65",x"69",x"69",x"89",x"89",x"89",x"a9",x"a9",x"a9",x"c5",x"c5",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"a4",x"a9",x"a9",x"a9",x"a9",x"89",x"89",x"89",x"89",x"69",x"69",x"6d",x"8d",x"8d",x"8d",x"8d",x"89",x"89",x"a9",x"a9",x"a9",x"c5",x"c5",x"c5",x"c0",x"c0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"84",x"a4",x"a8",x"a9",x"ad",x"ad",x"b2",x"b2",x"b2",x"d6",x"d6",x"db",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"d2",x"8d",x"04",x"20",x"80",x"a0",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"88",x"d0",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"ac",x"8c",x"88",x"68",x"68",x"68",x"44",x"44",x"44",x"44",x"40",x"40",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"44",x"88",x"b0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f5",x"d4",x"b0",x"8c",x"8c",x"8c",x"6c",x"68",x"68",x"48",x"44",x"40",x"20",x"20",x"20",x"20",x"68",x"ac",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"8c",x"8c",x"68",x"44",x"20",x"20",x"44",x"8c",x"b0",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f8",x"f9",x"f9",x"f9",x"f8",x"f4",x"f4",x"f4",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"b0",x"b0",x"90",x"8c",x"68",x"64",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"44",x"44",x"44",x"48",x"48",x"68",x"68",x"48",x"44",x"44",x"24",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"60",x"60",x"40",x"20",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"69",x"a9",x"a9",x"c9",x"c9",x"e5",x"e5",x"e5",x"e5",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"64",x"64",x"84",x"84",x"84",x"84",x"a4",x"a5",x"a5",x"a9",x"a9",x"a9",x"a9",x"a9",x"a9",x"a9",x"89",x"89",x"89",x"69",x"69",x"69",x"49",x"69",x"6d",x"8c",x"88",x"88",x"a8",x"a4",x"c4",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"88",x"89",x"b1",x"b2",x"b6",x"da",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"d2",x"8d",x"00",x"20",x"80",x"a0",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"88",x"cc",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"68",x"68",x"68",x"44",x"44",x"44",x"44",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"44",x"88",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"8c",x"8c",x"8c",x"6c",x"68",x"68",x"48",x"44",x"20",x"20",x"20",x"20",x"20",x"44",x"8c",x"b0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"b0",x"ac",x"8c",x"8c",x"8c",x"8c",x"68",x"68",x"20",x"20",x"44",x"8c",x"b0",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f8",x"f9",x"f9",x"f9",x"f9",x"f4",x"f4",x"f4",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"b0",x"b0",x"90",x"8c",x"8c",x"68",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"20",x"20",x"40",x"44",x"44",x"44",x"64",x"64",x"64",x"84",x"88",x"a9",x"a9",x"a9",x"c4",x"c4",x"e0",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"89",x"89",x"69",x"69",x"69",x"69",x"69",x"69",x"69",x"69",x"89",x"89",x"a9",x"a9",x"a9",x"a5",x"a4",x"a4",x"c4",x"c4",x"c4",x"c0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"84",x"84",x"89",x"a9",x"ad",x"cd",x"d2",x"d2",x"d6",x"d6",x"da",x"db",x"db",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"f6",x"8d",x"00",x"00",x"80",x"a0",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"80",x"80",x"80",x"84",x"ac",x"d0",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d0",x"b0",x"ac",x"8c",x"88",x"68",x"68",x"68",x"44",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"64",x"8c",x"d0",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"8c",x"8c",x"8c",x"6c",x"68",x"68",x"48",x"44",x"20",x"20",x"20",x"20",x"20",x"44",x"8c",x"b0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"b0",x"b0",x"ac",x"8c",x"8c",x"8c",x"8c",x"68",x"40",x"20",x"40",x"68",x"b0",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f8",x"f9",x"f9",x"f9",x"f9",x"f4",x"f4",x"f4",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"b0",x"b0",x"90",x"8c",x"8c",x"68",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"60",x"40",x"40",x"24",x"04",x"04",x"04",x"24",x"44",x"65",x"85",x"85",x"a5",x"c5",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"81",x"85",x"85",x"85",x"85",x"85",x"89",x"89",x"89",x"88",x"88",x"88",x"88",x"69",x"69",x"69",x"69",x"49",x"48",x"48",x"48",x"68",x"88",x"88",x"a8",x"c4",x"e4",x"e4",x"e4",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"64",x"64",x"64",x"68",x"89",x"8d",x"b2",x"d6",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"f6",x"ad",x"00",x"00",x"60",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"80",x"80",x"80",x"84",x"ac",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d0",x"d0",x"ac",x"8c",x"88",x"68",x"68",x"68",x"44",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"68",x"ac",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"8c",x"8c",x"8c",x"6c",x"68",x"68",x"48",x"44",x"20",x"20",x"20",x"20",x"20",x"40",x"68",x"ac",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"ac",x"ac",x"8c",x"8c",x"8c",x"68",x"44",x"20",x"20",x"44",x"8c",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f8",x"f9",x"f9",x"f9",x"f8",x"f4",x"f4",x"f4",x"f4",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"d0",x"b0",x"b0",x"90",x"8c",x"8c",x"68",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"20",x"20",x"20",x"24",x"44",x"44",x"44",x"44",x"64",x"64",x"85",x"85",x"84",x"a4",x"a4",x"c4",x"c4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"a4",x"a4",x"84",x"84",x"84",x"64",x"68",x"68",x"69",x"69",x"69",x"69",x"69",x"69",x"69",x"85",x"85",x"84",x"a4",x"a4",x"a4",x"c4",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"84",x"a8",x"a9",x"ad",x"b1",x"b2",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"f7",x"b2",x"00",x"00",x"60",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"84",x"a8",x"d0",x"d0",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"88",x"68",x"68",x"44",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"20",x"20",x"20",x"88",x"b0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"b0",x"ac",x"8c",x"8c",x"8c",x"68",x"68",x"68",x"44",x"44",x"20",x"20",x"20",x"20",x"20",x"20",x"64",x"8c",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f9",x"f8",x"f4",x"d4",x"f4",x"f8",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"ac",x"8c",x"8c",x"8c",x"8c",x"44",x"20",x"20",x"40",x"8c",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f8",x"f8",x"f9",x"f9",x"f9",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"b0",x"b0",x"90",x"8c",x"88",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"80",x"60",x"60",x"40",x"20",x"20",x"04",x"04",x"24",x"24",x"44",x"64",x"64",x"84",x"a4",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"84",x"84",x"84",x"64",x"68",x"84",x"84",x"84",x"84",x"84",x"68",x"68",x"68",x"68",x"68",x"69",x"69",x"69",x"89",x"89",x"85",x"a4",x"a4",x"c4",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"64",x"89",x"8d",x"b2",x"d6",x"da",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"fb",x"b2",x"20",x"00",x"40",x"60",x"80",x"80",x"60",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"84",x"a8",x"ac",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"88",x"68",x"64",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"8c",x"d0",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"6c",x"68",x"68",x"68",x"44",x"44",x"20",x"20",x"20",x"20",x"20",x"20",x"44",x"8c",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f9",x"f8",x"f4",x"f4",x"f4",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"b0",x"b0",x"ac",x"8c",x"8c",x"8c",x"8c",x"68",x"44",x"20",x"20",x"8c",x"b0",x"d4",x"d4",x"d4",x"d4",x"f4",x"f8",x"f8",x"f9",x"f9",x"f9",x"f8",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"b0",x"90",x"8c",x"88",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"a0",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"44",x"44",x"64",x"64",x"84",x"84",x"a4",x"a4",x"c4",x"c4",x"c0",x"c1",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"84",x"80",x"80",x"80",x"80",x"a0",x"a4",x"84",x"84",x"84",x"64",x"64",x"64",x"64",x"48",x"48",x"48",x"48",x"68",x"68",x"88",x"88",x"a4",x"a4",x"c4",x"c4",x"c4",x"c0",x"c0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"84",x"84",x"89",x"a9",x"ce",x"ce",x"d2",x"d6",x"d6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"fb",x"b2",x"20",x"00",x"40",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"88",x"ac",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"88",x"68",x"44",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"20",x"40",x"40",x"20",x"44",x"ac",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"8c",x"8c",x"8c",x"6c",x"68",x"68",x"48",x"44",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"68",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f9",x"f9",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"b0",x"b0",x"ac",x"8c",x"8c",x"8c",x"8c",x"68",x"44",x"20",x"20",x"68",x"b0",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f8",x"f9",x"f9",x"f9",x"f9",x"f8",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d0",x"b0",x"b0",x"b0",x"90",x"8c",x"88",x"44",x"20",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"20",x"20",x"00",x"00",x"04",x"24",x"44",x"44",x"64",x"84",x"84",x"a4",x"c4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"64",x"64",x"64",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"64",x"64",x"64",x"64",x"64",x"64",x"44",x"44",x"44",x"64",x"64",x"84",x"a4",x"a4",x"c4",x"c4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"60",x"64",x"64",x"68",x"89",x"8d",x"8d",x"b2",x"d6",x"f7",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"fb",x"b2",x"20",x"00",x"20",x"40",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"84",x"a8",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"ac",x"8c",x"68",x"68",x"44",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"68",x"b0",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"b0",x"8c",x"8c",x"8c",x"68",x"68",x"68",x"48",x"24",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"68",x"b0",x"d0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f9",x"f9",x"f8",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"68",x"68",x"20",x"20",x"68",x"8c",x"b0",x"d4",x"d4",x"d4",x"d4",x"f4",x"f8",x"f9",x"f9",x"f9",x"f9",x"f9",x"f4",x"f8",x"f8",x"f8",x"f9",x"f9",x"f4",x"d4",x"d0",x"b0",x"b0",x"b0",x"90",x"8c",x"68",x"44",x"20",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"60",x"60",x"40",x"20",x"00",x"00",x"00",x"00",x"04",x"24",x"24",x"24",x"44",x"64",x"64",x"84",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"84",x"84",x"84",x"84",x"84",x"64",x"64",x"44",x"44",x"24",x"24",x"24",x"44",x"44",x"64",x"84",x"84",x"a4",x"a4",x"a4",x"c0",x"c0",x"c0",x"c0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"60",x"60",x"60",x"80",x"80",x"80",x"84",x"a9",x"ad",x"ad",x"b2",x"b6",x"d6",x"d6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"b6",x"44",x"00",x"20",x"40",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"60",x"84",x"a8",x"cc",x"d0",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d0",x"d0",x"b0",x"ac",x"8c",x"88",x"68",x"68",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"64",x"8c",x"d0",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"8c",x"68",x"68",x"68",x"44",x"24",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"64",x"8c",x"b0",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f9",x"f9",x"f8",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"b0",x"b0",x"ac",x"8c",x"8c",x"8c",x"8c",x"68",x"20",x"20",x"44",x"8c",x"b0",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f9",x"f9",x"f9",x"f9",x"f9",x"f4",x"f4",x"f8",x"f8",x"f8",x"f9",x"f4",x"d4",x"b0",x"b0",x"b0",x"b0",x"90",x"8c",x"68",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"40",x"40",x"20",x"00",x"00",x"00",x"04",x"24",x"24",x"44",x"64",x"64",x"84",x"a4",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"84",x"84",x"84",x"84",x"84",x"64",x"64",x"64",x"64",x"44",x"44",x"44",x"44",x"44",x"44",x"64",x"84",x"a4",x"a4",x"c4",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"64",x"64",x"64",x"64",x"84",x"84",x"89",x"ad",x"b2",x"d6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"d6",x"44",x"20",x"20",x"40",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"60",x"84",x"88",x"ac",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d0",x"d0",x"b0",x"ac",x"8c",x"8c",x"68",x"68",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"64",x"88",x"b0",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"b0",x"ac",x"8c",x"8c",x"6c",x"68",x"68",x"68",x"44",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"44",x"8c",x"b0",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"f8",x"f9",x"f9",x"f8",x"f8",x"f4",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"68",x"44",x"20",x"44",x"68",x"b0",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f9",x"f9",x"f9",x"f9",x"f9",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"b0",x"90",x"8c",x"6c",x"48",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"60",x"60",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"80",x"60",x"40",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"60",x"84",x"80",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"84",x"84",x"64",x"64",x"44",x"44",x"24",x"24",x"24",x"24",x"44",x"64",x"84",x"a4",x"c4",x"c4",x"c0",x"c0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"84",x"89",x"ad",x"cd",x"d2",x"d6",x"d6",x"fb",x"fb",x"fb",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"d7",x"69",x"20",x"20",x"40",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"60",x"84",x"88",x"ac",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d0",x"d0",x"b0",x"ac",x"8c",x"8c",x"68",x"48",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"64",x"ac",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"8c",x"6c",x"68",x"68",x"68",x"44",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"44",x"68",x"b0",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f9",x"f9",x"f9",x"f8",x"f4",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"d4",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"68",x"44",x"20",x"20",x"44",x"b0",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f9",x"f9",x"f9",x"f9",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"b0",x"b0",x"b0",x"b0",x"90",x"8c",x"68",x"44",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"60",x"40",x"20",x"20",x"00",x"00",x"20",x"20",x"20",x"20",x"40",x"40",x"60",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"64",x"64",x"64",x"64",x"64",x"64",x"64",x"64",x"64",x"40",x"40",x"40",x"40",x"64",x"84",x"84",x"a4",x"c4",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"64",x"64",x"64",x"64",x"69",x"89",x"8d",x"b2",x"d6",x"fa",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"db",x"69",x"20",x"20",x"40",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"60",x"60",x"84",x"88",x"ac",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"d0",x"b0",x"ac",x"8c",x"6c",x"68",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"88",x"d0",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"d0",x"b0",x"ac",x"8c",x"8c",x"8c",x"6c",x"68",x"68",x"68",x"44",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"68",x"ac",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f9",x"f9",x"f9",x"f8",x"f4",x"f4",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"d4",x"b0",x"b0",x"8c",x"90",x"90",x"8c",x"6c",x"44",x"20",x"20",x"44",x"ac",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f9",x"f9",x"f9",x"f5",x"d4",x"d4",x"d4",x"d4",x"d4",x"d0",x"d0",x"b0",x"b0",x"b0",x"90",x"90",x"8c",x"68",x"44",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"20",x"20",x"00",x"00",x"00",x"00",x"20",x"20",x"40",x"60",x"60",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"64",x"64",x"64",x"40",x"40",x"40",x"44",x"44",x"44",x"44",x"44",x"60",x"80",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"60",x"40",x"40",x"60",x"60",x"80",x"84",x"89",x"8d",x"ad",x"b1",x"b2",x"d6",x"da",x"db",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"fb",x"8d",x"44",x"00",x"20",x"60",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"60",x"80",x"84",x"ac",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d0",x"d0",x"b0",x"b0",x"8c",x"6c",x"68",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"64",x"ac",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"d0",x"b0",x"ac",x"8c",x"8c",x"8c",x"6c",x"68",x"68",x"44",x"44",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"44",x"8c",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"f8",x"f9",x"f9",x"f9",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"b0",x"b0",x"b0",x"b0",x"90",x"8c",x"6c",x"44",x"20",x"20",x"20",x"8c",x"b0",x"b4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d5",x"f5",x"f5",x"d5",x"d4",x"d4",x"d0",x"d0",x"b0",x"b0",x"b0",x"b0",x"90",x"90",x"90",x"8c",x"6c",x"48",x"24",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"60",x"80",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"64",x"64",x"64",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"60",x"64",x"64",x"44",x"64",x"68",x"89",x"8d",x"ad",x"b2",x"d6",x"d6",x"db",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"fb",x"ce",x"65",x"00",x"00",x"60",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"60",x"84",x"a8",x"d0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"f9",x"f8",x"d4",x"d4",x"d4",x"d0",x"d0",x"b0",x"b0",x"8c",x"68",x"68",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"88",x"ac",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"8c",x"8c",x"68",x"68",x"68",x"44",x"40",x"20",x"20",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"68",x"b0",x"d4",x"d4",x"d4",x"f4",x"d4",x"d4",x"f8",x"f9",x"f9",x"f9",x"f5",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"d0",x"b0",x"b0",x"b0",x"b0",x"8c",x"6c",x"48",x"44",x"20",x"20",x"44",x"8c",x"b0",x"d4",x"d4",x"d0",x"b0",x"b0",x"d0",x"d4",x"d4",x"d4",x"d0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"8c",x"68",x"44",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"40",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"20",x"20",x"40",x"60",x"80",x"80",x"a0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"60",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"60",x"80",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"60",x"40",x"40",x"40",x"40",x"60",x"64",x"89",x"89",x"8d",x"b2",x"b2",x"d6",x"d6",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"f2",x"89",x"00",x"00",x"40",x"60",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"a8",x"b0",x"d0",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"fd",x"f9",x"f8",x"d4",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"8c",x"68",x"68",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"40",x"88",x"ac",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"d0",x"d0",x"b0",x"8c",x"8c",x"8c",x"8c",x"6c",x"68",x"68",x"44",x"44",x"20",x"20",x"20",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"68",x"b0",x"d0",x"d4",x"d4",x"f4",x"d4",x"d4",x"f8",x"f9",x"f9",x"f9",x"f5",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d0",x"b0",x"b0",x"b0",x"90",x"8c",x"6c",x"48",x"24",x"20",x"20",x"24",x"68",x"90",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"68",x"44",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"60",x"60",x"80",x"a0",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"84",x"64",x"64",x"64",x"69",x"69",x"89",x"8d",x"b2",x"b6",x"d6",x"db",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"f6",x"8d",x"20",x"00",x"40",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"88",x"ac",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"fd",x"fd",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"8c",x"8c",x"68",x"64",x"64",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"64",x"ac",x"f5",x"f9",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"6c",x"68",x"68",x"44",x"40",x"20",x"20",x"20",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"68",x"b0",x"d0",x"d4",x"d4",x"d4",x"d4",x"f4",x"f8",x"f9",x"f9",x"f9",x"f9",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f9",x"f9",x"d4",x"d0",x"b0",x"b0",x"b0",x"90",x"8c",x"6c",x"48",x"24",x"20",x"00",x"20",x"44",x"6c",x"90",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"90",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"6c",x"48",x"44",x"20",x"20",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"60",x"60",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"60",x"60",x"40",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"20",x"40",x"60",x"60",x"80",x"a0",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"80",x"80",x"80",x"60",x"60",x"40",x"20",x"20",x"20",x"20",x"24",x"20",x"40",x"60",x"80",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"a0",x"a0",x"80",x"80",x"60",x"40",x"40",x"40",x"40",x"60",x"84",x"a9",x"ad",x"cd",x"d2",x"d6",x"d7",x"fb",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"fb",x"b2",x"20",x"20",x"20",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"84",x"ac",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"f9",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"b0",x"ac",x"88",x"68",x"64",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"68",x"ac",x"d4",x"f9",x"f9",x"f9",x"f8",x"f8",x"f8",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"d0",x"d0",x"b0",x"ac",x"8c",x"8c",x"8c",x"8c",x"68",x"68",x"44",x"44",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"68",x"8c",x"b0",x"d4",x"d4",x"d4",x"d4",x"f4",x"f8",x"f9",x"f9",x"f9",x"f9",x"f9",x"f4",x"f4",x"f4",x"f8",x"f8",x"f9",x"f9",x"d5",x"b0",x"b0",x"b0",x"b0",x"8c",x"8c",x"6c",x"48",x"24",x"00",x"00",x"20",x"20",x"44",x"68",x"8c",x"b0",x"b0",x"b0",x"90",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"6c",x"48",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"a0",x"a0",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"60",x"60",x"80",x"80",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"84",x"64",x"68",x"69",x"69",x"6d",x"8d",x"b2",x"d2",x"f6",x"f6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"b6",x"40",x"20",x"20",x"40",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"84",x"88",x"ac",x"d0",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"d0",x"b0",x"8c",x"88",x"68",x"64",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"40",x"40",x"64",x"8c",x"d0",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"6c",x"68",x"68",x"44",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"44",x"8c",x"b0",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f9",x"f9",x"f9",x"f9",x"f9",x"f4",x"d4",x"d4",x"d4",x"f8",x"f9",x"f5",x"d5",x"b0",x"b0",x"b0",x"8c",x"8c",x"6c",x"68",x"44",x"20",x"00",x"00",x"00",x"20",x"20",x"44",x"68",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"6c",x"68",x"48",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"60",x"60",x"80",x"80",x"a0",x"c0",x"c0",x"a0",x"a0",x"80",x"60",x"40",x"40",x"20",x"00",x"00",x"00",x"00",x"20",x"20",x"40",x"40",x"60",x"80",x"a0",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"40",x"40",x"60",x"60",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"60",x"40",x"40",x"20",x"40",x"85",x"a9",x"89",x"ad",x"b2",x"b6",x"ba",x"db",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"d6",x"65",x"20",x"00",x"40",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"64",x"88",x"ac",x"d0",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"64",x"44",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"64",x"ac",x"d0",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"d4",x"b0",x"b0",x"ac",x"8c",x"8c",x"8c",x"8c",x"6c",x"68",x"44",x"24",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"44",x"68",x"b0",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f9",x"f9",x"f9",x"f9",x"f4",x"d4",x"d4",x"d4",x"d4",x"d5",x"d5",x"d0",x"b0",x"b0",x"b0",x"8c",x"8c",x"68",x"48",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"44",x"68",x"68",x"68",x"6c",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"6c",x"6c",x"68",x"48",x"44",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"40",x"40",x"40",x"60",x"80",x"80",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"84",x"84",x"84",x"89",x"69",x"69",x"69",x"8d",x"b2",x"d2",x"d6",x"d6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"db",x"a9",x"44",x"00",x"20",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"84",x"ac",x"d0",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"8c",x"88",x"64",x"64",x"44",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"64",x"88",x"ac",x"d0",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"d4",x"d0",x"b0",x"ac",x"8c",x"8c",x"8c",x"8c",x"6c",x"68",x"48",x"44",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"68",x"8c",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"f9",x"f9",x"f9",x"f9",x"f4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d0",x"b0",x"ac",x"b0",x"b0",x"8c",x"8c",x"68",x"44",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"44",x"44",x"48",x"68",x"68",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"68",x"68",x"48",x"24",x"20",x"20",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"40",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"40",x"40",x"60",x"80",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"40",x"60",x"80",x"a0",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"a0",x"80",x"60",x"60",x"60",x"40",x"40",x"64",x"89",x"8d",x"b2",x"d6",x"db",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"db",x"d2",x"69",x"00",x"20",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"a8",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f4",x"d4",x"d4",x"d0",x"b0",x"ac",x"ac",x"88",x"88",x"68",x"64",x"64",x"64",x"64",x"64",x"64",x"64",x"64",x"64",x"64",x"88",x"ac",x"d0",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"b0",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"68",x"44",x"24",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"44",x"8c",x"b0",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f9",x"f9",x"f9",x"d4",x"d4",x"d0",x"b0",x"b0",x"b0",x"b0",x"b0",x"ac",x"b0",x"b0",x"8c",x"8c",x"48",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"24",x"44",x"44",x"48",x"48",x"48",x"48",x"48",x"44",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"80",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a4",x"a4",x"a5",x"a9",x"89",x"89",x"8d",x"8d",x"92",x"b2",x"b6",x"d6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"d7",x"8d",x"00",x"00",x"40",x"60",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"a8",x"cc",x"d0",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d0",x"b0",x"ac",x"ac",x"ac",x"ac",x"ac",x"ac",x"ac",x"b0",x"b0",x"d0",x"d4",x"f4",x"f9",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"b0",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"68",x"48",x"44",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"20",x"20",x"68",x"b0",x"b4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"d4",x"d4",x"b0",x"b0",x"b0",x"b0",x"b0",x"ac",x"8c",x"8c",x"90",x"8c",x"8c",x"68",x"44",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"40",x"40",x"20",x"20",x"00",x"00",x"24",x"24",x"44",x"44",x"64",x"84",x"a4",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"40",x"20",x"20",x"20",x"40",x"40",x"60",x"60",x"80",x"a0",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"80",x"60",x"60",x"40",x"40",x"40",x"64",x"69",x"89",x"ad",x"b2",x"d6",x"d7",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"b2",x"20",x"00",x"20",x"40",x"60",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"84",x"ac",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d0",x"b0",x"b0",x"ac",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"68",x"44",x"24",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"20",x"44",x"8c",x"b0",x"b4",x"d4",x"d4",x"d4",x"b0",x"b0",x"d4",x"d4",x"d4",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"8c",x"8c",x"90",x"8c",x"8c",x"68",x"68",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"a0",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"a0",x"a4",x"84",x"88",x"89",x"89",x"8d",x"8d",x"b2",x"b6",x"d6",x"db",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"b6",x"40",x"20",x"20",x"40",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"84",x"a8",x"d0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"b0",x"b0",x"ac",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"68",x"48",x"24",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"20",x"44",x"68",x"8c",x"b0",x"b0",x"b4",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"90",x"90",x"90",x"90",x"8c",x"8c",x"8c",x"90",x"8c",x"68",x"48",x"44",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"60",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"60",x"80",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"40",x"60",x"80",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"40",x"60",x"64",x"88",x"ad",x"ad",x"d2",x"d6",x"d6",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"d6",x"69",x"20",x"00",x"20",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"84",x"a8",x"b0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"d0",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"68",x"48",x"44",x"20",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"20",x"44",x"68",x"6c",x"8c",x"b0",x"b0",x"b0",x"90",x"90",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"68",x"44",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"44",x"40",x"60",x"60",x"60",x"80",x"80",x"a0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"84",x"88",x"89",x"ad",x"ad",x"ae",x"b2",x"b2",x"d6",x"d6",x"fb",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"ae",x"44",x"00",x"20",x"40",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"84",x"88",x"ac",x"d0",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d0",x"b0",x"b0",x"ac",x"8c",x"8c",x"8c",x"8c",x"6c",x"68",x"68",x"44",x"24",x"20",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"48",x"68",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"68",x"48",x"44",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"80",x"60",x"40",x"40",x"20",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"44",x"64",x"84",x"84",x"a4",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"40",x"60",x"80",x"80",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"60",x"60",x"60",x"64",x"64",x"69",x"8d",x"b2",x"d6",x"f6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"d6",x"89",x"20",x"20",x"40",x"60",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"88",x"ac",x"d0",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"b0",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"68",x"48",x"44",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"44",x"68",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"6c",x"6c",x"6c",x"68",x"48",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"64",x"64",x"64",x"84",x"84",x"84",x"a4",x"a4",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"84",x"84",x"89",x"a9",x"ad",x"ad",x"b2",x"b2",x"b6",x"d6",x"d7",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"ad",x"20",x"20",x"40",x"60",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"ac",x"d0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"fd",x"f9",x"f9",x"f9",x"f9",x"f8",x"f4",x"d4",x"d4",x"d0",x"b0",x"b0",x"ac",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"68",x"44",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"44",x"68",x"68",x"68",x"6c",x"8c",x"8c",x"8c",x"6c",x"6c",x"68",x"68",x"68",x"48",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"80",x"80",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"60",x"40",x"40",x"20",x"24",x"04",x"04",x"04",x"24",x"44",x"44",x"64",x"84",x"a4",x"c4",x"c4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"80",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"64",x"64",x"64",x"68",x"8d",x"8d",x"b2",x"d6",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"b6",x"44",x"20",x"20",x"40",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"60",x"84",x"ac",x"d0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"f9",x"f9",x"f8",x"d4",x"d4",x"d0",x"b0",x"b0",x"ac",x"8c",x"8c",x"8c",x"8c",x"6c",x"68",x"68",x"44",x"24",x"20",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"44",x"48",x"68",x"68",x"68",x"68",x"68",x"44",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"a0",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"44",x"44",x"44",x"44",x"44",x"64",x"64",x"64",x"64",x"84",x"84",x"84",x"a4",x"a4",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"80",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"84",x"89",x"a9",x"ad",x"b2",x"d2",x"d2",x"d6",x"d6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"6d",x"24",x"20",x"40",x"60",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"60",x"60",x"60",x"88",x"b0",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"fd",x"fd",x"f9",x"f9",x"d4",x"d4",x"b0",x"b0",x"b0",x"ac",x"8c",x"8c",x"8c",x"8c",x"6c",x"68",x"48",x"44",x"24",x"20",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"44",x"44",x"44",x"44",x"44",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"60",x"60",x"40",x"40",x"24",x"24",x"24",x"24",x"24",x"48",x"48",x"64",x"84",x"a4",x"a4",x"c4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"a0",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"60",x"60",x"60",x"60",x"64",x"64",x"89",x"89",x"ad",x"b2",x"d6",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"48",x"20",x"20",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"88",x"ac",x"d0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"ff",x"ff",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"d4",x"d4",x"b0",x"b0",x"b0",x"b0",x"b0",x"8c",x"8c",x"8c",x"6c",x"6c",x"48",x"44",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"20",x"24",x"24",x"24",x"44",x"44",x"44",x"64",x"68",x"68",x"89",x"89",x"a5",x"a4",x"c4",x"c4",x"c4",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"40",x"60",x"60",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"84",x"84",x"89",x"ad",x"b2",x"b2",x"d2",x"d6",x"d6",x"db",x"db",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"d6",x"6d",x"20",x"40",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"84",x"a8",x"d0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fe",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"fd",x"f9",x"f9",x"f9",x"d4",x"d4",x"b0",x"b0",x"ac",x"ac",x"b0",x"8c",x"8c",x"8c",x"6c",x"6c",x"68",x"48",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"40",x"24",x"24",x"24",x"05",x"09",x"29",x"48",x"68",x"88",x"88",x"a9",x"c9",x"c5",x"e5",x"e5",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"40",x"20",x"20",x"20",x"40",x"40",x"60",x"80",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"60",x"60",x"60",x"64",x"64",x"89",x"8d",x"b1",x"b2",x"d6",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"b2",x"44",x"40",x"40",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"84",x"88",x"b0",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"fd",x"fd",x"f9",x"f9",x"f9",x"d5",x"d4",x"d4",x"b0",x"b0",x"ac",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"68",x"48",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"80",x"80",x"80",x"a0",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"20",x"24",x"24",x"44",x"44",x"44",x"44",x"68",x"69",x"69",x"89",x"89",x"89",x"89",x"a9",x"a8",x"c8",x"c8",x"c4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"40",x"20",x"20",x"40",x"40",x"60",x"60",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"80",x"80",x"60",x"60",x"60",x"80",x"a0",x"a0",x"a4",x"a9",x"ad",x"ad",x"b2",x"b2",x"b6",x"d6",x"da",x"db",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"d6",x"89",x"64",x"40",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"88",x"ac",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"fd",x"fd",x"fd",x"f9",x"f9",x"d9",x"d9",x"d4",x"b0",x"b0",x"b0",x"ac",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"68",x"48",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"44",x"24",x"28",x"29",x"49",x"49",x"69",x"69",x"89",x"a9",x"a9",x"c9",x"c9",x"e9",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"20",x"20",x"20",x"40",x"40",x"60",x"80",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"60",x"60",x"44",x"44",x"64",x"84",x"a5",x"a9",x"ad",x"b2",x"d6",x"db",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"b2",x"89",x"40",x"40",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"88",x"ac",x"d0",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fc",x"fc",x"fc",x"f8",x"fc",x"fc",x"fc",x"fd",x"fd",x"fd",x"fc",x"fc",x"fc",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"fd",x"fd",x"fd",x"fd",x"f9",x"d9",x"d5",x"b4",x"b0",x"b0",x"b0",x"ac",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"68",x"44",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"a0",x"a0",x"80",x"80",x"60",x"40",x"20",x"24",x"24",x"24",x"28",x"29",x"49",x"49",x"49",x"6d",x"8d",x"8d",x"ad",x"a9",x"a9",x"c9",x"c5",x"c4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"20",x"00",x"00",x"00",x"40",x"60",x"60",x"60",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"84",x"89",x"ad",x"b1",x"b2",x"b6",x"d6",x"db",x"db",x"db",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"ad",x"60",x"40",x"40",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"ac",x"d0",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"d9",x"d5",x"b4",x"b0",x"b0",x"b0",x"ac",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"68",x"44",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"80",x"80",x"64",x"44",x"24",x"28",x"28",x"28",x"49",x"4d",x"6d",x"6d",x"8d",x"ad",x"cd",x"e9",x"e9",x"e9",x"e8",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"40",x"40",x"20",x"20",x"20",x"60",x"80",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"84",x"84",x"64",x"64",x"64",x"64",x"64",x"89",x"8d",x"b2",x"d6",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"d6",x"89",x"40",x"40",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"a8",x"ac",x"d0",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"fd",x"fd",x"fd",x"fd",x"fd",x"fd",x"f9",x"f9",x"f9",x"f5",x"d5",x"d4",x"b0",x"b0",x"b0",x"b0",x"ac",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"48",x"44",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"60",x"60",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"44",x"24",x"24",x"24",x"49",x"69",x"69",x"69",x"69",x"8d",x"8d",x"8d",x"ad",x"ad",x"c9",x"c9",x"c9",x"c4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"40",x"60",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"60",x"60",x"40",x"40",x"60",x"60",x"60",x"84",x"88",x"ad",x"ad",x"b2",x"b6",x"d6",x"da",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"b2",x"64",x"20",x"40",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"a8",x"ac",x"d0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fd",x"fd",x"fd",x"fd",x"fd",x"f9",x"f9",x"f9",x"d5",x"d4",x"b0",x"b0",x"b0",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"68",x"48",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"64",x"64",x"65",x"49",x"49",x"29",x"49",x"69",x"8d",x"8d",x"8d",x"ad",x"ad",x"cd",x"ed",x"e9",x"e9",x"e9",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"64",x"64",x"44",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"80",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"80",x"80",x"64",x"44",x"44",x"44",x"64",x"69",x"89",x"8d",x"b2",x"d6",x"da",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"f6",x"89",x"40",x"40",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"60",x"80",x"88",x"ac",x"d0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"fd",x"fd",x"fd",x"fd",x"f9",x"f9",x"f9",x"d5",x"d5",x"b0",x"b0",x"b0",x"b0",x"ac",x"ac",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"48",x"44",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"40",x"40",x"60",x"60",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"60",x"40",x"20",x"44",x"44",x"48",x"49",x"49",x"6d",x"6d",x"8d",x"8d",x"ad",x"cd",x"ce",x"ce",x"ed",x"ed",x"ed",x"e9",x"e9",x"e5",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"64",x"64",x"84",x"84",x"80",x"80",x"80",x"80",x"81",x"80",x"80",x"60",x"40",x"40",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"80",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"80",x"60",x"40",x"20",x"40",x"60",x"84",x"89",x"ad",x"ae",x"d2",x"d2",x"d6",x"d7",x"fb",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"b2",x"64",x"40",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"84",x"ac",x"d0",x"d4",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"d9",x"d5",x"d5",x"b4",x"b0",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"68",x"48",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"40",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"84",x"64",x"45",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"8d",x"ad",x"ad",x"cd",x"ed",x"e9",x"e9",x"e9",x"e9",x"e9",x"e8",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"60",x"80",x"80",x"80",x"80",x"84",x"84",x"84",x"84",x"64",x"64",x"64",x"64",x"60",x"64",x"64",x"64",x"60",x"60",x"60",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"a0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"84",x"84",x"64",x"44",x"44",x"68",x"69",x"ad",x"b2",x"d6",x"fb",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"d6",x"8d",x"64",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"a8",x"d0",x"d4",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"f9",x"d9",x"d5",x"d5",x"b4",x"b0",x"b0",x"b0",x"90",x"90",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"6c",x"68",x"48",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"60",x"80",x"a0",x"a0",x"c0",x"c0",x"a0",x"a0",x"80",x"60",x"40",x"40",x"24",x"24",x"28",x"49",x"4d",x"6d",x"6d",x"6e",x"b2",x"b2",x"b2",x"d2",x"d2",x"ce",x"ee",x"ed",x"e9",x"e9",x"e9",x"e5",x"e5",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"40",x"40",x"24",x"24",x"44",x"44",x"60",x"80",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"80",x"60",x"40",x"40",x"40",x"40",x"60",x"84",x"89",x"ad",x"ce",x"d2",x"d6",x"db",x"db",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"d6",x"8d",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"60",x"84",x"88",x"b0",x"d4",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f4",x"f4",x"f4",x"f5",x"f5",x"f5",x"d5",x"d5",x"d5",x"d4",x"d4",x"d4",x"d4",x"d4",x"b0",x"b0",x"b0",x"90",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"68",x"68",x"48",x"44",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"a0",x"84",x"84",x"84",x"64",x"68",x"49",x"49",x"4d",x"6d",x"6d",x"92",x"92",x"92",x"b2",x"d2",x"ed",x"ed",x"ed",x"ed",x"e9",x"e9",x"e9",x"e5",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"e0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"84",x"84",x"84",x"68",x"69",x"69",x"89",x"8d",x"ae",x"d2",x"d6",x"f7",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"d2",x"84",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"60",x"60",x"84",x"ac",x"b0",x"b4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f8",x"f8",x"f8",x"f4",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"d4",x"d4",x"d4",x"d4",x"d4",x"d0",x"d0",x"d0",x"d0",x"d4",x"d4",x"d4",x"d4",x"d4",x"d4",x"b4",x"b0",x"b0",x"b0",x"b0",x"b0",x"ac",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"6c",x"68",x"44",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"80",x"80",x"80",x"a0",x"a0",x"80",x"80",x"60",x"60",x"40",x"40",x"24",x"24",x"49",x"4d",x"4d",x"6d",x"92",x"92",x"b2",x"d2",x"d2",x"d2",x"f2",x"ee",x"ee",x"ed",x"ed",x"e9",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"64",x"64",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"80",x"80",x"80",x"84",x"84",x"84",x"64",x"64",x"64",x"64",x"64",x"84",x"84",x"84",x"80",x"a0",x"a0",x"a0",x"c0",x"c0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"40",x"40",x"60",x"85",x"89",x"ad",x"b2",x"d6",x"f6",x"fb",x"fb",x"fb",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"b1",x"64",x"40",x"60",x"60",x"80",x"80",x"80",x"80",x"60",x"84",x"ac",x"b0",x"b4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f8",x"f8",x"f4",x"d4",x"b4",x"b0",x"b0",x"90",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"90",x"90",x"90",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"6c",x"68",x"48",x"48",x"44",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"84",x"84",x"64",x"64",x"69",x"69",x"69",x"6d",x"6d",x"6d",x"92",x"92",x"b2",x"b2",x"d2",x"f2",x"ee",x"ed",x"ed",x"e9",x"e9",x"e9",x"e9",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"84",x"64",x"64",x"64",x"64",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"a4",x"a4",x"a4",x"a4",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"84",x"84",x"84",x"89",x"89",x"89",x"89",x"8d",x"b2",x"b6",x"d6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"8d",x"44",x"60",x"60",x"60",x"80",x"80",x"80",x"60",x"84",x"88",x"b0",x"d4",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"f9",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"b0",x"b0",x"8c",x"8c",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"ac",x"ac",x"ac",x"ac",x"ac",x"ac",x"ac",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"68",x"48",x"44",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"40",x"44",x"44",x"49",x"4d",x"4d",x"71",x"72",x"92",x"b2",x"b6",x"d6",x"d2",x"f2",x"f2",x"f2",x"ed",x"ed",x"e9",x"e9",x"e5",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"80",x"80",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"a4",x"a0",x"c4",x"c4",x"e4",x"e4",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"40",x"40",x"40",x"40",x"40",x"64",x"69",x"8d",x"b2",x"d2",x"d6",x"fb",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"b6",x"8d",x"60",x"40",x"60",x"80",x"80",x"80",x"60",x"80",x"88",x"b0",x"d4",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f9",x"f4",x"d4",x"b0",x"b0",x"8c",x"8c",x"6c",x"6c",x"6c",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"68",x"68",x"68",x"48",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"80",x"80",x"84",x"84",x"84",x"85",x"89",x"89",x"89",x"8d",x"8d",x"92",x"92",x"92",x"b2",x"b2",x"d2",x"d2",x"f2",x"f2",x"ed",x"ed",x"ed",x"e9",x"e9",x"e5",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"85",x"88",x"88",x"88",x"84",x"84",x"84",x"84",x"a4",x"a4",x"a4",x"a4",x"c4",x"c4",x"c4",x"c4",x"c4",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"84",x"84",x"89",x"89",x"89",x"8d",x"8d",x"b2",x"b2",x"b6",x"db",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"d6",x"64",x"40",x"60",x"80",x"80",x"60",x"60",x"60",x"88",x"ac",x"b0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f9",x"f8",x"f4",x"d4",x"b0",x"b0",x"8c",x"8c",x"6c",x"68",x"68",x"6c",x"6c",x"8c",x"8c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"8c",x"8c",x"8c",x"8c",x"8c",x"8c",x"6c",x"6c",x"6c",x"6c",x"68",x"48",x"44",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"40",x"40",x"40",x"60",x"60",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"65",x"69",x"69",x"6d",x"6e",x"92",x"b6",x"b6",x"b6",x"d6",x"f6",x"f6",x"f2",x"f2",x"f2",x"ee",x"ed",x"e9",x"e9",x"e9",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"64",x"84",x"84",x"85",x"85",x"85",x"85",x"85",x"85",x"85",x"89",x"89",x"89",x"89",x"89",x"88",x"88",x"88",x"a4",x"a4",x"a4",x"c4",x"c4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"64",x"88",x"89",x"8d",x"b1",x"d6",x"f6",x"f6",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"b2",x"89",x"60",x"60",x"60",x"60",x"60",x"80",x"84",x"ac",x"b0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"d4",x"b0",x"b0",x"8c",x"8c",x"6c",x"68",x"68",x"6c",x"8c",x"6c",x"68",x"68",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"48",x"44",x"44",x"44",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"80",x"84",x"84",x"84",x"84",x"88",x"89",x"89",x"8d",x"8d",x"8e",x"92",x"92",x"92",x"b2",x"b2",x"d2",x"d2",x"f2",x"f2",x"ed",x"ed",x"ed",x"e9",x"e9",x"e9",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"85",x"85",x"85",x"85",x"89",x"89",x"89",x"89",x"89",x"89",x"a9",x"a9",x"a9",x"a9",x"a9",x"a9",x"c4",x"c4",x"c4",x"c4",x"c4",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"a0",x"a0",x"a4",x"a4",x"a5",x"a9",x"a9",x"ad",x"ad",x"b2",x"b6",x"b6",x"b6",x"da",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"64",x"20",x"60",x"60",x"80",x"80",x"84",x"88",x"b0",x"d0",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"d4",x"d4",x"b0",x"90",x"8c",x"8c",x"8c",x"6c",x"6c",x"6c",x"68",x"64",x"64",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"68",x"48",x"44",x"44",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"44",x"44",x"48",x"69",x"6d",x"71",x"91",x"96",x"b6",x"b6",x"d6",x"d6",x"f6",x"f6",x"f6",x"f2",x"f2",x"ed",x"ed",x"e9",x"e9",x"e5",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"84",x"84",x"84",x"84",x"84",x"84",x"85",x"85",x"89",x"89",x"89",x"a5",x"a5",x"a5",x"a9",x"a9",x"a9",x"a9",x"a9",x"a9",x"a9",x"a8",x"a4",x"a4",x"c4",x"c4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"84",x"85",x"a9",x"ce",x"d2",x"d6",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"ad",x"64",x"40",x"40",x"60",x"80",x"60",x"88",x"ac",x"d0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"d4",x"d4",x"b0",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"6c",x"84",x"80",x"60",x"60",x"64",x"64",x"44",x"44",x"44",x"44",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"64",x"64",x"65",x"69",x"89",x"89",x"8d",x"8d",x"92",x"92",x"92",x"b2",x"b6",x"b6",x"b6",x"d6",x"d6",x"f2",x"f2",x"ed",x"ed",x"e9",x"e9",x"e5",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a4",x"a4",x"a4",x"84",x"a4",x"a4",x"a5",x"85",x"85",x"85",x"89",x"89",x"89",x"89",x"89",x"89",x"89",x"89",x"89",x"89",x"89",x"a9",x"a9",x"a9",x"a9",x"c9",x"c9",x"c9",x"c4",x"c4",x"c4",x"c4",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"84",x"84",x"89",x"89",x"a9",x"ad",x"ad",x"b2",x"b2",x"d6",x"d6",x"db",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"b1",x"44",x"40",x"60",x"60",x"60",x"84",x"ac",x"d0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"d4",x"b0",x"b0",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"84",x"80",x"80",x"80",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"20",x"20",x"20",x"20",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"60",x"64",x"44",x"48",x"49",x"4d",x"6d",x"72",x"92",x"b2",x"b6",x"d6",x"f7",x"f7",x"f7",x"d6",x"d6",x"d2",x"d2",x"f1",x"ed",x"e9",x"e5",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a4",x"a4",x"84",x"84",x"84",x"84",x"85",x"85",x"a5",x"a9",x"a9",x"89",x"89",x"89",x"89",x"89",x"ad",x"ad",x"ad",x"ad",x"8d",x"8d",x"8d",x"8d",x"88",x"a8",x"a8",x"a8",x"c8",x"c8",x"e4",x"e4",x"e4",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"80",x"60",x"80",x"80",x"80",x"60",x"64",x"64",x"88",x"89",x"ad",x"b2",x"d6",x"d6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"da",x"ad",x"64",x"60",x"40",x"60",x"84",x"ac",x"d0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"d4",x"b0",x"b0",x"90",x"8c",x"8c",x"8c",x"8c",x"84",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"64",x"64",x"64",x"89",x"89",x"89",x"8d",x"8d",x"92",x"92",x"96",x"b6",x"b6",x"d2",x"d2",x"d2",x"f2",x"f2",x"ee",x"ee",x"ee",x"e9",x"e9",x"e9",x"e9",x"e5",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a4",x"a4",x"a4",x"84",x"84",x"89",x"89",x"89",x"89",x"89",x"89",x"a9",x"a9",x"ad",x"ad",x"8d",x"8d",x"8d",x"8d",x"ad",x"ad",x"a9",x"c9",x"c9",x"c9",x"c9",x"c9",x"c9",x"c4",x"e4",x"e4",x"c4",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"a0",x"a0",x"80",x"84",x"84",x"89",x"a9",x"ad",x"b1",x"b2",x"b2",x"d6",x"d6",x"da",x"db",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"f6",x"ad",x"60",x"40",x"40",x"64",x"ac",x"b0",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"f9",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"8c",x"68",x"64",x"60",x"60",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"60",x"60",x"40",x"40",x"40",x"60",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"40",x"60",x"60",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"80",x"84",x"64",x"48",x"49",x"49",x"4d",x"6e",x"72",x"92",x"96",x"b6",x"da",x"fa",x"fa",x"f6",x"f6",x"f2",x"ed",x"ed",x"e9",x"e9",x"e5",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"84",x"84",x"84",x"84",x"84",x"84",x"a5",x"a5",x"85",x"89",x"89",x"89",x"89",x"89",x"89",x"8d",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"c9",x"c9",x"c9",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"60",x"60",x"60",x"60",x"60",x"64",x"84",x"84",x"89",x"ad",x"b2",x"b2",x"d6",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"f7",x"ae",x"85",x"40",x"40",x"68",x"ac",x"b0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"f9",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"d4",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"8c",x"48",x"24",x"24",x"20",x"20",x"40",x"40",x"40",x"60",x"60",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"64",x"64",x"64",x"69",x"89",x"8d",x"8d",x"92",x"92",x"b2",x"b2",x"b2",x"b2",x"d2",x"d2",x"d2",x"f2",x"f2",x"ee",x"ed",x"e9",x"e9",x"e9",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a4",x"a4",x"84",x"84",x"85",x"85",x"85",x"89",x"89",x"89",x"89",x"89",x"89",x"89",x"89",x"8d",x"8d",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"c9",x"c9",x"c9",x"c9",x"e9",x"e9",x"e5",x"e5",x"e4",x"e0",x"e0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"84",x"89",x"89",x"ad",x"ae",x"b2",x"d2",x"d6",x"d6",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"f7",x"ae",x"64",x"40",x"64",x"88",x"b0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"f9",x"f9",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"d4",x"d4",x"b0",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"48",x"28",x"24",x"04",x"04",x"00",x"00",x"00",x"20",x"40",x"40",x"60",x"80",x"80",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"60",x"64",x"65",x"69",x"69",x"6d",x"71",x"92",x"96",x"b6",x"d6",x"d6",x"f6",x"f6",x"f2",x"f2",x"f2",x"ed",x"ed",x"e9",x"e5",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"84",x"84",x"84",x"84",x"84",x"89",x"89",x"89",x"89",x"89",x"89",x"89",x"89",x"89",x"8d",x"8d",x"8d",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"cd",x"cd",x"c9",x"c9",x"c9",x"c9",x"c9",x"e4",x"e5",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"a0",x"80",x"60",x"60",x"40",x"40",x"60",x"64",x"84",x"89",x"ad",x"d2",x"d2",x"d6",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"b2",x"89",x"44",x"68",x"b0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"fd",x"f9",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"d4",x"b0",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"8d",x"69",x"69",x"69",x"49",x"49",x"49",x"44",x"44",x"44",x"44",x"44",x"40",x"40",x"40",x"40",x"40",x"40",x"44",x"44",x"44",x"44",x"44",x"44",x"64",x"64",x"68",x"89",x"89",x"8d",x"8d",x"8e",x"8e",x"b2",x"b2",x"b2",x"b2",x"d6",x"d2",x"d2",x"f2",x"f2",x"ed",x"ed",x"ed",x"e9",x"e8",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a4",x"a4",x"a4",x"a4",x"84",x"84",x"88",x"89",x"89",x"89",x"89",x"89",x"8d",x"8d",x"8d",x"8d",x"8d",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"cd",x"cd",x"cd",x"c9",x"e9",x"e9",x"e9",x"e5",x"e5",x"e5",x"e4",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"84",x"84",x"88",x"89",x"ad",x"b2",x"b2",x"b2",x"d6",x"d6",x"db",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"b2",x"68",x"68",x"b0",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"fd",x"f9",x"f9",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"f4",x"d4",x"d4",x"d4",x"b0",x"b0",x"90",x"8c",x"8c",x"ac",x"cd",x"cd",x"ad",x"ad",x"ad",x"8d",x"8d",x"6d",x"6d",x"69",x"49",x"49",x"49",x"49",x"29",x"29",x"29",x"29",x"29",x"49",x"49",x"49",x"49",x"49",x"4d",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"d6",x"d6",x"d6",x"f6",x"f6",x"f2",x"f2",x"f2",x"ed",x"e9",x"e9",x"e5",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"84",x"84",x"84",x"84",x"84",x"a4",x"a4",x"a9",x"a9",x"a9",x"a9",x"a9",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"b1",x"ad",x"ad",x"cd",x"cd",x"cd",x"cd",x"c9",x"e9",x"e9",x"e5",x"e5",x"e5",x"e4",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"80",x"60",x"40",x"40",x"40",x"40",x"64",x"89",x"8d",x"ad",x"d2",x"d2",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"b1",x"b0",x"d0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"f9",x"f9",x"f9",x"f9",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"d4",x"b0",x"b0",x"90",x"8c",x"6c",x"8c",x"a8",x"ac",x"cd",x"cd",x"cd",x"ce",x"d2",x"d2",x"d2",x"b2",x"b2",x"b2",x"92",x"96",x"96",x"b6",x"b6",x"96",x"96",x"96",x"96",x"b6",x"b6",x"b6",x"b6",x"b6",x"d6",x"d6",x"d6",x"d6",x"f2",x"f2",x"ed",x"ed",x"ed",x"e9",x"e9",x"e5",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a4",x"a4",x"a4",x"a4",x"84",x"84",x"89",x"89",x"89",x"89",x"89",x"a9",x"a9",x"a9",x"a9",x"ad",x"ad",x"ad",x"ad",x"ad",x"ae",x"b2",x"b2",x"d1",x"cd",x"cd",x"cd",x"ed",x"ed",x"ed",x"e9",x"e5",x"e5",x"e5",x"e4",x"e4",x"e4",x"e0",x"c0",x"c0",x"a0",x"80",x"80",x"60",x"60",x"60",x"80",x"80",x"84",x"84",x"89",x"8d",x"ad",x"b2",x"d2",x"d6",x"d6",x"db",x"fb",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"da",x"b0",x"b0",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"fd",x"fd",x"f9",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"f4",x"d4",x"d4",x"b0",x"b0",x"90",x"8c",x"6c",x"88",x"88",x"a8",x"c8",x"e9",x"ed",x"ed",x"ed",x"ed",x"ee",x"f2",x"f2",x"f6",x"f6",x"d6",x"fb",x"fa",x"f6",x"f6",x"f6",x"f6",x"f6",x"f6",x"f6",x"f6",x"f6",x"f6",x"f2",x"f2",x"f2",x"ed",x"ed",x"e9",x"e9",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a4",x"84",x"84",x"84",x"89",x"89",x"89",x"89",x"89",x"89",x"89",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"b2",x"d2",x"d2",x"d2",x"cd",x"cd",x"cd",x"ed",x"e9",x"e9",x"e9",x"e5",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"80",x"60",x"60",x"40",x"40",x"44",x"84",x"a9",x"ad",x"ad",x"d2",x"d6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fa",x"d5",x"b4",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"fd",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f4",x"d4",x"d4",x"b4",x"b0",x"90",x"90",x"8c",x"8c",x"88",x"a8",x"c8",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e8",x"e9",x"e9",x"e9",x"ed",x"ed",x"ed",x"ed",x"ed",x"ed",x"ed",x"ed",x"ed",x"e9",x"e9",x"e9",x"e9",x"e9",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a4",x"a4",x"84",x"84",x"84",x"84",x"84",x"84",x"89",x"89",x"a9",x"a9",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"b1",x"b1",x"b1",x"b1",x"b1",x"b1",x"d1",x"d1",x"ed",x"ed",x"ed",x"ed",x"e9",x"e9",x"e9",x"e5",x"e4",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"60",x"60",x"60",x"60",x"60",x"60",x"84",x"84",x"a9",x"ad",x"ae",x"b2",x"b2",x"d2",x"d6",x"fb",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"d6",x"b5",x"b4",x"d4",x"d8",x"f8",x"f4",x"f4",x"f4",x"f9",x"f9",x"fd",x"fd",x"fd",x"fc",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f4",x"d4",x"d4",x"b4",x"b0",x"b0",x"90",x"8c",x"6c",x"6c",x"88",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"84",x"84",x"84",x"84",x"84",x"88",x"68",x"68",x"89",x"89",x"89",x"a9",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"cd",x"cd",x"cd",x"d1",x"d1",x"d1",x"d1",x"d1",x"cd",x"ad",x"ad",x"cd",x"ed",x"e9",x"e9",x"e9",x"e8",x"e4",x"c4",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"40",x"40",x"40",x"40",x"44",x"64",x"69",x"8d",x"ae",x"d2",x"d6",x"fb",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"da",x"d5",x"b4",x"d4",x"d4",x"f8",x"f4",x"f4",x"f8",x"f9",x"f9",x"fd",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f4",x"d4",x"d4",x"b4",x"b0",x"b0",x"90",x"8c",x"90",x"90",x"8c",x"a8",x"c4",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"84",x"84",x"84",x"84",x"84",x"a5",x"a5",x"a5",x"a9",x"a9",x"a9",x"a9",x"ad",x"ad",x"ad",x"ad",x"ad",x"cd",x"cd",x"d1",x"d1",x"b1",x"b1",x"b1",x"b1",x"b1",x"d1",x"d1",x"d1",x"ed",x"ed",x"e9",x"e9",x"e5",x"e5",x"e4",x"e0",x"e0",x"c0",x"a0",x"a0",x"80",x"60",x"60",x"40",x"40",x"40",x"40",x"60",x"84",x"a9",x"8d",x"ad",x"b2",x"d2",x"d6",x"d6",x"db",x"db",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fa",x"d5",x"b4",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f9",x"f9",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f9",x"f8",x"d4",x"d4",x"b4",x"b0",x"b0",x"90",x"8c",x"90",x"90",x"8c",x"88",x"a4",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"84",x"84",x"84",x"84",x"84",x"84",x"88",x"88",x"89",x"a9",x"a9",x"a9",x"a9",x"ad",x"ad",x"ad",x"ad",x"cd",x"cd",x"d2",x"d2",x"d2",x"d2",x"d2",x"d1",x"d1",x"d1",x"cd",x"cd",x"cd",x"cd",x"cd",x"c9",x"c9",x"e9",x"e5",x"e0",x"e0",x"e0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"64",x"44",x"44",x"44",x"44",x"64",x"89",x"ad",x"d2",x"d6",x"da",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d5",x"b0",x"b4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f9",x"f9",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"f8",x"d4",x"d4",x"d4",x"b0",x"b0",x"90",x"8c",x"8c",x"8c",x"88",x"88",x"84",x"80",x"a0",x"a0",x"c0",x"c0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"84",x"84",x"84",x"84",x"89",x"89",x"89",x"89",x"a9",x"a9",x"a9",x"a9",x"ad",x"ad",x"ad",x"ad",x"ad",x"ae",x"d2",x"d2",x"d2",x"d2",x"d1",x"d1",x"d1",x"d1",x"cd",x"ed",x"e9",x"e9",x"e9",x"e5",x"e5",x"e5",x"e4",x"c0",x"c0",x"a0",x"a0",x"80",x"60",x"60",x"40",x"40",x"40",x"60",x"60",x"85",x"ad",x"ce",x"d2",x"d6",x"d6",x"d6",x"da",x"db",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"da",x"b0",x"b4",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fd",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f9",x"f8",x"f4",x"d4",x"d4",x"b0",x"b0",x"90",x"8c",x"8c",x"8c",x"88",x"88",x"84",x"84",x"80",x"80",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"e0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a4",x"a4",x"a4",x"a4",x"84",x"84",x"84",x"84",x"84",x"89",x"89",x"89",x"89",x"8d",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"b2",x"b2",x"ae",x"cd",x"cd",x"cd",x"cd",x"cd",x"ed",x"ed",x"cd",x"cd",x"cd",x"c9",x"c9",x"e5",x"e4",x"e4",x"e0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"64",x"64",x"44",x"44",x"69",x"69",x"8d",x"b2",x"f6",x"f7",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"da",x"b5",x"b4",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"fd",x"fd",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"b0",x"b0",x"b0",x"8c",x"90",x"90",x"8c",x"68",x"68",x"88",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"80",x"80",x"a4",x"a4",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"a9",x"a9",x"a9",x"a9",x"a9",x"a9",x"ad",x"ad",x"ad",x"ad",x"ad",x"b1",x"b2",x"b2",x"b2",x"d2",x"d1",x"d1",x"cd",x"cd",x"ed",x"ed",x"ed",x"e9",x"e9",x"e9",x"e4",x"e4",x"e0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"60",x"60",x"60",x"40",x"60",x"64",x"84",x"a9",x"cd",x"d2",x"f2",x"d6",x"db",x"db",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fa",x"b5",x"b4",x"d4",x"d4",x"d4",x"f8",x"f8",x"f8",x"f8",x"f9",x"f9",x"fd",x"fd",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"b0",x"b0",x"b0",x"90",x"90",x"6c",x"6c",x"68",x"68",x"88",x"88",x"85",x"84",x"84",x"84",x"84",x"84",x"64",x"64",x"64",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"84",x"88",x"88",x"89",x"89",x"89",x"89",x"a9",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"cd",x"cd",x"d1",x"d1",x"d1",x"cd",x"cd",x"cd",x"cd",x"ed",x"ed",x"e9",x"e9",x"e9",x"e4",x"e4",x"e4",x"c4",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"84",x"84",x"64",x"68",x"69",x"69",x"8d",x"b1",x"d6",x"f6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"b5",x"b4",x"b4",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f8",x"f9",x"fd",x"fe",x"fd",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"b0",x"b0",x"b0",x"90",x"8c",x"6c",x"6c",x"68",x"68",x"88",x"89",x"a5",x"a5",x"a5",x"89",x"89",x"89",x"69",x"68",x"68",x"89",x"a9",x"89",x"89",x"89",x"89",x"a9",x"a9",x"a9",x"a9",x"a9",x"ad",x"ad",x"ad",x"ad",x"ad",x"8d",x"ad",x"b1",x"b1",x"b1",x"b1",x"d1",x"d1",x"cd",x"ed",x"ed",x"e9",x"e9",x"e9",x"e5",x"e4",x"e4",x"e4",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"64",x"89",x"ad",x"ad",x"d2",x"f6",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"df",x"df",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"d6",x"b5",x"b4",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f9",x"fd",x"fe",x"fd",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"b0",x"b0",x"b0",x"90",x"8c",x"6c",x"68",x"68",x"68",x"88",x"a9",x"a9",x"a9",x"a9",x"a9",x"89",x"89",x"89",x"89",x"89",x"89",x"89",x"89",x"89",x"89",x"a9",x"a9",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"b1",x"b1",x"b1",x"cd",x"cd",x"cd",x"cd",x"e9",x"e9",x"e9",x"e5",x"c5",x"c4",x"c4",x"c4",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"84",x"84",x"85",x"89",x"89",x"89",x"8d",x"b1",x"b2",x"d6",x"da",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"da",x"d5",x"b4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f9",x"f9",x"fe",x"fd",x"fd",x"f9",x"f8",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d0",x"b0",x"b0",x"b0",x"90",x"8c",x"6c",x"6c",x"68",x"68",x"84",x"a9",x"a9",x"a9",x"a9",x"a9",x"a9",x"a9",x"a9",x"a9",x"a9",x"8d",x"8d",x"8d",x"8d",x"8d",x"8d",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"ad",x"d1",x"d1",x"cd",x"ed",x"e9",x"e5",x"e4",x"e0",x"e0",x"c0",x"c0",x"a0",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"64",x"64",x"89",x"ad",x"ae",x"d2",x"d6",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fa",x"d5",x"b4",x"d4",x"d4",x"d4",x"f4",x"f4",x"f8",x"f8",x"f8",x"f9",x"fe",x"fd",x"fd",x"f9",x"f8",x"f8",x"f8",x"f8",x"f4",x"d4",x"d4",x"b0",x"b0",x"b0",x"90",x"8c",x"6c",x"6c",x"68",x"84",x"84",x"a4",x"c4",x"c5",x"c5",x"c5",x"c4",x"c4",x"c4",x"c4",x"c5",x"c9",x"c9",x"c9",x"c9",x"c9",x"c9",x"c9",x"c9",x"c9",x"c9",x"c9",x"c9",x"c9",x"c9",x"c9",x"c9",x"c9",x"e9",x"e9",x"e4",x"c4",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"80",x"80",x"80",x"84",x"84",x"68",x"89",x"89",x"8d",x"8d",x"b2",x"b2",x"d6",x"db",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"da",x"b4",x"b4",x"d4",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f9",x"fe",x"fd",x"fd",x"f9",x"f8",x"d4",x"d4",x"d4",x"d4",x"d4",x"d0",x"b0",x"b0",x"90",x"90",x"8c",x"6c",x"68",x"64",x"84",x"a0",x"c0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e0",x"e4",x"e4",x"e4",x"e5",x"e5",x"e5",x"e5",x"e5",x"e5",x"e5",x"e5",x"e5",x"e5",x"e5",x"e4",x"e4",x"e4",x"e4",x"e4",x"e0",x"e0",x"c0",x"a0",x"a0",x"80",x"80",x"60",x"60",x"60",x"84",x"84",x"a9",x"a9",x"a9",x"d2",x"d6",x"d6",x"f7",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"da",x"b0",x"b4",x"d4",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f9",x"fe",x"fe",x"fd",x"f9",x"d8",x"d4",x"d4",x"d4",x"d4",x"d4",x"b0",x"b0",x"90",x"8c",x"8c",x"8c",x"68",x"48",x"64",x"a4",x"c4",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"c0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"a0",x"80",x"84",x"84",x"84",x"89",x"8d",x"ad",x"b1",x"b2",x"d2",x"d6",x"d6",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"da",x"b4",x"b4",x"d4",x"d4",x"d4",x"f4",x"f8",x"f8",x"f8",x"f9",x"f9",x"fd",x"fd",x"f9",x"d8",x"d4",x"d4",x"d4",x"d4",x"d4",x"b0",x"b0",x"8c",x"8c",x"8c",x"8c",x"6c",x"48",x"68",x"ad",x"a9",x"a4",x"80",x"80",x"60",x"60",x"60",x"60",x"80",x"80",x"a0",x"a0",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"80",x"60",x"60",x"60",x"60",x"60",x"64",x"64",x"89",x"8d",x"b1",x"b6",x"d6",x"db",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fa",x"d5",x"b4",x"b4",x"b4",x"d4",x"d4",x"f4",x"f8",x"f8",x"f9",x"f9",x"f9",x"f9",x"f9",x"d4",x"d4",x"d4",x"b4",x"b0",x"b0",x"b0",x"90",x"8c",x"8c",x"6c",x"68",x"6c",x"91",x"b6",x"d6",x"d2",x"d2",x"ad",x"ad",x"8d",x"8d",x"8d",x"8d",x"89",x"89",x"a9",x"a4",x"84",x"84",x"84",x"84",x"88",x"88",x"88",x"89",x"89",x"89",x"89",x"a9",x"a9",x"a9",x"ad",x"ad",x"b2",x"b2",x"b6",x"d6",x"db",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"da",x"b5",x"b0",x"b0",x"b0",x"b4",x"d4",x"d4",x"d4",x"d4",x"d4",x"d5",x"d5",x"d4",x"d4",x"d0",x"b0",x"b0",x"b0",x"90",x"90",x"90",x"90",x"8c",x"68",x"68",x"b6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"db",x"d6",x"d6",x"b2",x"b2",x"b2",x"b2",x"b2",x"b2",x"b2",x"b2",x"b2",x"b2",x"d6",x"d6",x"d6",x"d6",x"f7",x"fb",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fe",x"d5",x"b0",x"90",x"90",x"b0",x"b4",x"d4",x"d4",x"d4",x"d0",x"d0",x"d0",x"d0",x"b0",x"b0",x"b0",x"b0",x"90",x"8c",x"8c",x"6c",x"6c",x"8c",x"91",x"b1",x"da",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"fb",x"fb",x"fb",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"da",x"b5",x"90",x"90",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"b0",x"90",x"90",x"8c",x"8c",x"6c",x"6c",x"8c",x"b1",x"d6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"b1",x"8d",x"8c",x"8c",x"8c",x"8c",x"b0",x"b0",x"b0",x"90",x"b0",x"90",x"8c",x"8c",x"6c",x"6c",x"6c",x"8c",x"b1",x"b6",x"da",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"d6",x"b1",x"8c",x"68",x"6c",x"8c",x"8c",x"90",x"8c",x"8c",x"90",x"8c",x"8c",x"6c",x"68",x"6c",x"8d",x"b5",x"da",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"b1",x"8c",x"8c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"6c",x"8c",x"91",x"b5",x"da",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"da",x"b5",x"91",x"8c",x"6c",x"6c",x"6c",x"6c",x"6c",x"8d",x"91",x"d6",x"fb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"fb",x"da",x"d6",x"b6",x"d6",x"da",x"da",x"da",x"da",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff")
);

constant object : object_form := (
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111100000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111110000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111001111111111100000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111000111111111100000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111100111111111110000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111100111111111110000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111100111111111110000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111100111111111110000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111110011111111111000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111000000111111111111111111110011111111111000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111101111111111111111111111011111111111100000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111001111111111100000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111001111111111100000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111001111111111100000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111101111111111110000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000001111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100000111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111110000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000011111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111111111111111111111110001100000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111111111111111111111111111111111111111111111111111111111111111001100000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100"),
("000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100"),
("000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100"),
("000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100"),
("000000000000000000000000000000000000000000000000000000000000000000001111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("000000000000000000000000000000000000000000000000000000000000001111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("000000000000000000000000000000000000000000000000000000001111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000"),
("000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000"),
("000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000"),
("000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000"),
("000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000"),
("000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000"),
("000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000"),
("000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000"),
("000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000"),
("000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000"),
("000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000"),
("000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000"),
("000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000"),
("000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000"),
("000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000"),
("000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000"),
("000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000"),
("000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000"),
("000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000"),
("000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000"),
("000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100010000000000"),
("000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000"),
("000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000"),
("000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000"),
("000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000"),
("000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000"),
("000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000"),
("000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000"),
("000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000"),
("000000000000111111111111111111111111111111111111111111111110000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000"),
("000000000001111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000"),
("000000000001111111111111111111111111111111111111111110000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000"),
("000000000011111111111111111111111111111111111111111100000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000"),
("000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000"),
("000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000"),
("000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000"),
("000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000"),
("000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000"),
("000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000"),
("000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000"),
("000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000"),
("000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000"),
("000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000"),
("000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000"),
("000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000"),
("000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000"),
("000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000"),
("000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000"),
("000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000"),
("000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000"),
("000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000"),
("001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000"),
("001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000"),
("001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000"),
("011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000"),
("011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000"),
("011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000"),
("011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000"),
("011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000"),
("011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000"),
("011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000010000000000000000000000000000000000000000000000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000011111111111111111111111111111111111111111111111111111111111110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000111000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000001111111111111111111111111110000000011111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000001111111111111111111111111110000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000")
);

signal bCoord_X : integer := 0;-- offset from start position 
signal bCoord_Y : integer := 0;

signal drawing_X : std_logic := '0';
signal drawing_Y : std_logic := '0';
	
signal objectEndX : integer;
signal objectEndY : integer;

begin

-- Calculate object end boundaries
objectEndX	<= object_X_size+ObjectStartX;
objectEndY	<= object_Y_size+ObjectStartY;

-- Signals drawing_X[Y] are active when obects coordinates are being crossed

-- test if ooCoord is in the rectangle defined by Start and End 
	drawing_X	<= '1' when  (oCoord_X  >= ObjectStartX) and  (oCoord_X < objectEndX) else '0';
    drawing_Y	<= '1' when  (oCoord_Y  >= ObjectStartY) and  (oCoord_Y < objectEndY) else '0';

-- calculate offset from start corner 
	bCoord_X 	<= (oCoord_X - ObjectStartX) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 
	bCoord_Y 	<= (oCoord_Y - ObjectStartY) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 


process ( RESETn, CLK)

  		
   begin
	if RESETn = '0' then
	    mVGA_RGB	<=  (others => '0') ; 	
		drawing_request	<=  '0' ;

		elsif rising_edge(CLK) then
			mVGA_RGB	<=  object_colors(bCoord_Y , bCoord_X);	--get from colors table 
			drawing_request	<= object(bCoord_Y , bCoord_X) and drawing_X and drawing_Y ; -- get from mask table if inside rectangle  
	end if;

  end process;

		
end behav;
