module controller 	(
			input	wire 	ENABLE,
			input	wire	reset,
			input	wire	fifo_Empty,
			input	wire	fifo_full,
			input 	wire	ps2_done,
			input 	wire	ps2_error,
			output	wire	DONE,
			output	wire	read,
			output	wire	write
			);



endmodule
