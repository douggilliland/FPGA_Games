--------------------------------------
-- SinTable.vhd
-- Written by Gadi and Eran Tuchman.
-- All rights reserved, Copyright 2009
--------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all ;

entity sintable is
port(
  CLK     					: in std_logic;
  resetN 					: in std_logic;
  ADDR    					: in std_logic_vector(7 downto 0);
  Q       					: out std_logic_vector(15 downto 0)
);
end sintable;

architecture arch of sintable is
constant array_size 			: integer := 256 ;

type table_type is array(0 to array_size - 1) of std_logic_vector(15 downto 0);
signal sin_table				: table_type;
signal Q_tmp       			:  std_logic_vector(15 downto 0) ;



begin
 
   
  sintable_proc: process(resetN, CLK)
    constant sin_table : table_type := (
X"C180",
X"C2F7",
X"C469",
X"C5D4",
X"C739",
X"C899",
X"C9F3",
X"CB47",
X"CC96",
X"CDDF",
X"CF22",
X"D060",
X"D199",
X"D2CC",
X"D3FA",
X"D523",
X"D646",
X"D764",
X"D87D",
X"D991",
X"DAA0",
X"DBA9",
X"DCAE",
X"DDAE",
X"DEA9",
X"DF9F",
X"E091",
X"E17D",
X"E265",
X"E349",
X"E428",
X"E502",
X"E5D8",
X"E6A9",
X"E776",
X"E83E",
X"E902",
X"E9C2",
X"EA7E",
X"EB35",
X"EBE9",
X"EC98",
X"ED44",
X"EDEB",
X"EE8E",
X"EF2E",
X"EFC9",
X"F061",
X"F0F5",
X"F186",
X"F213",
X"F29C",
X"F321",
X"F3A3",
X"F422",
X"F49D",
X"F515",
X"F589",
X"F5FB",
X"F668",
X"F6D3",
X"F73B",
X"F79F",
X"F801",
X"F85F",
X"F8BB",
X"F914",
X"F969",
X"F9BC",
X"FA0C",
X"FA5A",
X"FAA5",
X"FAED",
X"FB33",
X"FB76",
X"FBB6",
X"FBF4",
X"FC30",
X"FC6A",
X"FCA1",
X"FCD6",
X"FD08",
X"FD39",
X"FD67",
X"FD93",
X"FDBE",
X"FDE6",
X"FE0D",
X"FE31",
X"FE54",
X"FE75",
X"FE94",
X"FEB2",
X"FECD",
X"FEE8",
X"FF01",
X"FF18",
X"FF2E",
X"FF42",
X"FF55",
X"FF67",
X"FF77",
X"FF86",
X"FF95",
X"FFA1",
X"FFAD",
X"FFB8",
X"FFC2",
X"FFCB",
X"FFD3",
X"FFDA",
X"FFE1",
X"FFE6",
X"FFEB",
X"FFEF",
X"FFF3",
X"FFF6",
X"FFF9",
X"FFFB",
X"FFFD",
X"FFFE",
X"FFFF",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0001",
X"0002",
X"0003",
X"0005",
X"0007",
X"000A",
X"000D",
X"0011",
X"0015",
X"001A",
X"001F",
X"0026",
X"002D",
X"0035",
X"003E",
X"0048",
X"0053",
X"005F",
X"006B",
X"007A",
X"0089",
X"0099",
X"00AB",
X"00BE",
X"00D2",
X"00E8",
X"00FF",
X"0118",
X"0133",
X"014E",
X"016C",
X"018B",
X"01AC",
X"01CF",
X"01F3",
X"021A",
X"0242",
X"026D",
X"0299",
X"02C7",
X"02F8",
X"032A",
X"035F",
X"0396",
X"03D0",
X"040C",
X"044A",
X"048A",
X"04CD",
X"0513",
X"055B",
X"05A6",
X"05F4",
X"0644",
X"0697",
X"06EC",
X"0745",
X"07A1",
X"07FF",
X"0861",
X"08C5",
X"092D",
X"0998",
X"0A05",
X"0A77",
X"0AEB",
X"0B63",
X"0BDE",
X"0C5D",
X"0CDF",
X"0D64",
X"0DED",
X"0E7A",
X"0F0B",
X"0F9F",
X"1037",
X"10D2",
X"1172",
X"1215",
X"12BC",
X"1368",
X"1417",
X"14CB",
X"1582",
X"163E",
X"16FE",
X"17C2",
X"188A",
X"1957",
X"1A28",
X"1AFE",
X"1BD8",
X"1CB7",
X"1D9B",
X"1E83",
X"1F6F",
X"2061",
X"2157",
X"2252",
X"2352",
X"2457",
X"2560",
X"266F",
X"2783",
X"289C",
X"29BA",
X"2ADD",
X"2C06",
X"2D34",
X"2E67",
X"2FA0",
X"30DE",
X"3221",
X"336A",
X"34B9",
X"360D",
X"3767",
X"38C7",
X"3A2C",
X"3B97",
X"3D09",
X"3E80",
X"3FFC");

 
 begin

    if (resetN='0') then
		Q_tmp <= ( others => '0');
    elsif(rising_edge(CLK)) then
--      if (ENA='1') then
		Q_tmp <= sin_table(conv_integer(ADDR));
--      end if;
   end if;
  end process;
 Q <= Q_tmp; 

		   
end arch;