library IEEE;
use IEEE.STD_LOGIC_1164.all;
--use IEEE.std_logic_unsigned.all;
--use ieee.numeric_std.all;
--use ieee.std_logic_arith.all;
-- Alex Grinshpun April 2017
-- Dudy Nov 13 2017


entity score  is
port 	(
		--////////////////////	Clock Input	 	////////////////////	
	   	CLK  		: in std_logic;
		RESETn		: in std_logic;
		oCoord_X	: in integer;
		oCoord_Y	: in integer;
		ObjectStartX   : in integer ;
	   ObjectStartY	: in integer ; 
	   digit   : in integer ; 	
		drawing_request	: out std_logic ;
		mVGA_RGB 	: out std_logic_vector(7 downto 0)

		
	); 
end score ;

architecture behav of score is 



constant ObjectStartY : integer := 10;

constant object_X_size : integer := 20;
constant object_Y_size : integer := 15;

--one heart

type ram_array0 is array(0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic_vector(7 downto 0);
constant object_colors0: ram_array0 := ( 
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"64",x"a4",x"c4",x"a4",x"a4",x"a4",x"a4",x"84",x"84",x"84",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"a4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"64",x"64",x"a4",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"20",x"20",x"60",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"a4",x"20",x"e8",x"e8",x"64",x"00",x"00"),
(x"00",x"00",x"00",x"c8",x"c4",x"40",x"00",x"40",x"64",x"64",x"64",x"64",x"60",x"20",x"c4",x"e8",x"e8",x"a4",x"00",x"00"),
(x"00",x"00",x"00",x"e8",x"e8",x"e8",x"a4",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"e8",x"e8",x"e8",x"a4",x"00",x"00"),
(x"00",x"00",x"00",x"e8",x"e8",x"e8",x"c4",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"e8",x"e8",x"e8",x"84",x"00",x"00"),
(x"00",x"00",x"20",x"e8",x"e8",x"e8",x"a4",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"e8",x"e8",x"e8",x"84",x"00",x"00"),
(x"00",x"00",x"20",x"e8",x"e8",x"e8",x"a4",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"e8",x"e8",x"e8",x"84",x"00",x"00"),
(x"00",x"00",x"40",x"e8",x"e8",x"e8",x"84",x"00",x"00",x"00",x"00",x"00",x"00",x"60",x"e8",x"e8",x"e8",x"64",x"00",x"00"),
(x"00",x"00",x"40",x"e8",x"e8",x"e8",x"84",x"00",x"00",x"00",x"00",x"00",x"00",x"64",x"e8",x"e8",x"e8",x"60",x"00",x"00"),
(x"00",x"00",x"60",x"e8",x"e8",x"e8",x"64",x"00",x"00",x"00",x"00",x"00",x"00",x"64",x"e8",x"e8",x"e8",x"40",x"00",x"00"),
(x"00",x"00",x"64",x"e8",x"e8",x"e8",x"60",x"00",x"00",x"00",x"00",x"00",x"00",x"84",x"e8",x"e8",x"e8",x"40",x"00",x"00"),
(x"00",x"00",x"84",x"e8",x"e8",x"a4",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"c4",x"e8",x"e8",x"40",x"00",x"00"),
(x"00",x"00",x"40",x"a4",x"40",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"84",x"c4",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"40",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00"),
(x"00",x"00",x"64",x"e8",x"e8",x"84",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"84",x"c4",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"84",x"e8",x"e8",x"e8",x"40",x"00",x"00",x"00",x"00",x"00",x"00",x"c4",x"e8",x"e8",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"84",x"e8",x"e8",x"e8",x"40",x"00",x"00",x"00",x"00",x"00",x"00",x"c4",x"e8",x"e8",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"84",x"e8",x"e8",x"e8",x"40",x"00",x"00",x"00",x"00",x"00",x"00",x"c4",x"e8",x"e8",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"84",x"e8",x"e8",x"e8",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"c8",x"e8",x"e8",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"a4",x"e8",x"e8",x"e8",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"e8",x"e8",x"e8",x"e8",x"00",x"00",x"00"),
(x"00",x"00",x"a4",x"e8",x"e8",x"e8",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"e8",x"e8",x"e8",x"e8",x"00",x"00",x"00"),
(x"00",x"00",x"a4",x"e8",x"e8",x"e8",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"e8",x"e8",x"e8",x"e8",x"00",x"00",x"00"),
(x"00",x"00",x"a4",x"e8",x"e8",x"e8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"e8",x"e8",x"e8",x"c4",x"00",x"00",x"00"),
(x"00",x"00",x"a4",x"e8",x"a4",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"c4",x"e8",x"e8",x"c4",x"00",x"00",x"00"),
(x"00",x"00",x"64",x"40",x"20",x"a4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"84",x"40",x"e8",x"e8",x"84",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"84",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"40",x"a4",x"c8",x"20",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"20",x"84",x"a4",x"a4",x"a4",x"a4",x"c4",x"c4",x"c4",x"c4",x"84",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00")


);


type object_form0 is array (0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic;
constant object0 : object_form0 := (
("00000000000000000000"),
("00000000000000000000"),
("00000111111111100000"),
("00001111111111111000"),
("00011111111111111100"),
("00011101111111111100"),
("00011110000001111100"),
("00011110000001111100"),
("00111110000001111100"),
("00111110000001111100"),
("00111110000001111100"),
("00111110000001111100"),
("00111110000001111100"),
("00111110000001111100"),
("00111100000001111100"),
("00111000000000011100"),
("00000000000000000000"),
("00010000000000001000"),
("00111100000001111100"),
("00111110000001111100"),
("00111110000001111100"),
("00111110000001111100"),
("00111110000001111100"),
("00111110000001111000"),
("00111110000001111000"),
("00111110000001111000"),
("00111100000001111000"),
("00111111111101111000"),
("00111111111111111000"),
("00011111111111111000"),
("00011111111111000000"),
("00000000000000000000"),
("00000000000000000000")
);

type ram_array1 is array(0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic_vector(7 downto 0);  

-- 8 bit - color definition : "RRRGGGBB"  
constant object_colors1: ram_array1 := ( 
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"64",x"a4",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"e8",x"e8",x"64",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"c4",x"e8",x"e8",x"a4",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"e8",x"e8",x"e8",x"a4",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"e8",x"e8",x"e8",x"84",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"e8",x"e8",x"e8",x"84",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"e8",x"e8",x"e8",x"84",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"60",x"e8",x"e8",x"e8",x"64",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"64",x"e8",x"e8",x"e8",x"60",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"64",x"e8",x"e8",x"e8",x"40",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"84",x"e8",x"e8",x"e8",x"40",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"c4",x"e8",x"e8",x"40",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"84",x"c4",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"84",x"c4",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"c4",x"e8",x"e8",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"c4",x"e8",x"e8",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"c4",x"e8",x"e8",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"c8",x"e8",x"e8",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"e8",x"e8",x"e8",x"e8",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"e8",x"e8",x"e8",x"e8",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"e8",x"e8",x"e8",x"e8",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"e8",x"e8",x"e8",x"c4",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"c4",x"e8",x"e8",x"c4",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"e8",x"e8",x"84",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"a4",x"c8",x"20",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00")


);


-- one bit mask  0 - off 1 dispaly 
type object_form1 is array (0 to object1_Y_size - 1 , 0 to object1_X_size - 1) of std_logic;
constant object1 : object_form1 := (
("00000000000000000000"),
("00000000000000000000"),
("00000000000000000000"),
("00000000000000011000"),
("00000000000000111100"),
("00000000000000111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000000011100"),
("00000000000000000000"),
("00000000000000001000"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111000"),
("00000000000001111000"),
("00000000000001111000"),
("00000000000001111000"),
("00000000000001111000"),
("00000000000001111000"),
("00000000000000111000"),
("00000000000000000000"),
("00000000000000000000"),
("00000000000000000000")

);

----two hears
type ram_array2 is array(0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic_vector(7 downto 0);

constant object_colors2: ram_array2 := ( 
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"64",x"a4",x"c4",x"a4",x"a4",x"a4",x"a4",x"84",x"84",x"84",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"a4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"64",x"64",x"a4",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"64",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"a4",x"20",x"e8",x"e8",x"64",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"64",x"64",x"64",x"64",x"60",x"20",x"c4",x"e8",x"e8",x"a4",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"e8",x"e8",x"e8",x"a4",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"e8",x"e8",x"e8",x"84",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"e8",x"e8",x"e8",x"84",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"e8",x"e8",x"e8",x"84",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"60",x"e8",x"e8",x"e8",x"64",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"64",x"e8",x"e8",x"e8",x"60",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"64",x"e8",x"e8",x"e8",x"40",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"84",x"e8",x"e8",x"e8",x"40",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"c4",x"e8",x"e8",x"40",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"20",x"c4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"84",x"20",x"64",x"c4",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"60",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"40",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"40",x"20",x"40",x"c4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"84",x"20",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"64",x"e8",x"e8",x"64",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"84",x"e8",x"e8",x"e8",x"40",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"84",x"e8",x"e8",x"e8",x"40",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"84",x"e8",x"e8",x"e8",x"40",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"84",x"e8",x"e8",x"e8",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"a4",x"e8",x"e8",x"e8",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"a4",x"e8",x"e8",x"e8",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"a4",x"e8",x"e8",x"e8",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"a4",x"e8",x"e8",x"e8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"a4",x"e8",x"a4",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"64",x"40",x"20",x"a4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"84",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"84",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"40",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"20",x"84",x"a4",x"a4",x"a4",x"a4",x"c4",x"c4",x"c4",x"c4",x"84",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00")


);


-- one bit mask  0 - off 1 dispaly 
type object_form2 is array (0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic;
constant object2 : object_form2 := (
("00000000000000000000"),
("00000000000000000000"),
("00000111111111100000"),
("00001111111111111000"),
("00000111111111111100"),
("00000001111111111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000001111111111100"),
("00000111111111111100"),
("00001111111111110000"),
("00011111111111110000"),
("00111100011110000000"),
("00111110000000000000"),
("00111110000000000000"),
("00111110000000000000"),
("00111110000000000000"),
("00111110000000000000"),
("00111110000000000000"),
("00111110000000000000"),
("00111100000000000000"),
("00111111111100000000"),
("00111111111110000000"),
("00011111111111000000"),
("00011111111111000000"),
("00000000000000000000"),
("00000000000000000000")
     

);

------3 hearts
type ram_array3 is array(0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic_vector(7 downto 0);
constant object_colors3: ram_array3 := ( 
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"64",x"a4",x"c4",x"a4",x"a4",x"a4",x"a4",x"84",x"84",x"84",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"a4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"64",x"64",x"a4",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"64",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"a4",x"20",x"e8",x"e8",x"64",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"64",x"64",x"64",x"64",x"60",x"20",x"c4",x"e8",x"e8",x"a4",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"e8",x"e8",x"e8",x"a4",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"e8",x"e8",x"e8",x"84",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"e8",x"e8",x"e8",x"84",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"e8",x"e8",x"e8",x"84",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"60",x"e8",x"e8",x"e8",x"64",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"64",x"e8",x"e8",x"e8",x"60",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"64",x"e8",x"e8",x"e8",x"40",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"84",x"e8",x"e8",x"e8",x"40",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"c4",x"e8",x"e8",x"40",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"20",x"c4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"84",x"20",x"64",x"c4",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"60",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"40",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"40",x"c4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"84",x"20",x"20",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"64",x"c4",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"c4",x"e8",x"e8",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"c4",x"e8",x"e8",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"c4",x"e8",x"e8",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"c8",x"e8",x"e8",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"e8",x"e8",x"e8",x"e8",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"e8",x"e8",x"e8",x"e8",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"e8",x"e8",x"e8",x"e8",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"e8",x"e8",x"e8",x"c4",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"c4",x"e8",x"e8",x"c4",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"20",x"a4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"84",x"40",x"e8",x"e8",x"84",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"a4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"40",x"a4",x"c8",x"20",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"20",x"84",x"a4",x"a4",x"a4",x"a4",x"c4",x"c4",x"c4",x"c4",x"84",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00")



);


type object_form3 is array (0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic;
constant object3 : object_form3 := (
("00000000000000000000"),
("00000000000000000000"),
("00000111111111100000"),
("00001111111111111000"),
("00000111111111111100"),
("00000001111111111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000001111111111100"),
("00000111111111111100"),
("00001111111111110000"),
("00000111111111111000"),
("00000000011111111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111000"),
("00000000000001111000"),
("00000000000001111000"),
("00000000000001111000"),
("00000011111101111000"),
("00001111111111111000"),
("00011111111111111000"),
("00011111111111000000"),
("00000000000000000000"),
("00000000000000000000")

);

type ram_array4 is array(0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic_vector(7 downto 0);
constant object_colors4: ram_array4 := ( 

(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"64",x"a4",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"e8",x"e8",x"64",x"00",x"00"),
(x"00",x"00",x"00",x"c8",x"c4",x"60",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"c4",x"e8",x"e8",x"a4",x"00",x"00"),
(x"00",x"00",x"00",x"e8",x"e8",x"e8",x"a4",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"e8",x"e8",x"e8",x"a4",x"00",x"00"),
(x"00",x"00",x"00",x"e8",x"e8",x"e8",x"c4",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"e8",x"e8",x"e8",x"84",x"00",x"00"),
(x"00",x"00",x"20",x"e8",x"e8",x"e8",x"a4",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"e8",x"e8",x"e8",x"84",x"00",x"00"),
(x"00",x"00",x"20",x"e8",x"e8",x"e8",x"a4",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"e8",x"e8",x"e8",x"84",x"00",x"00"),
(x"00",x"00",x"40",x"e8",x"e8",x"e8",x"84",x"00",x"00",x"00",x"00",x"00",x"00",x"60",x"e8",x"e8",x"e8",x"64",x"00",x"00"),
(x"00",x"00",x"40",x"e8",x"e8",x"e8",x"84",x"00",x"00",x"00",x"00",x"00",x"00",x"64",x"e8",x"e8",x"e8",x"60",x"00",x"00"),
(x"00",x"00",x"60",x"e8",x"e8",x"e8",x"64",x"00",x"00",x"00",x"00",x"00",x"00",x"64",x"e8",x"e8",x"e8",x"40",x"00",x"00"),
(x"00",x"00",x"64",x"e8",x"e8",x"e8",x"60",x"00",x"00",x"00",x"00",x"00",x"00",x"84",x"e8",x"e8",x"e8",x"40",x"00",x"00"),
(x"00",x"00",x"84",x"e8",x"e8",x"a4",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"c4",x"e8",x"e8",x"40",x"00",x"00"),
(x"00",x"00",x"40",x"a4",x"40",x"20",x"a4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"84",x"20",x"64",x"c4",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"60",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"40",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"40",x"c4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"84",x"20",x"20",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"64",x"c4",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"c4",x"e8",x"e8",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"c4",x"e8",x"e8",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"c4",x"e8",x"e8",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"c8",x"e8",x"e8",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"e8",x"e8",x"e8",x"e8",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"e8",x"e8",x"e8",x"e8",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"e8",x"e8",x"e8",x"e8",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"e8",x"e8",x"e8",x"c4",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"c4",x"e8",x"e8",x"c4",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"e8",x"e8",x"84",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"a4",x"c8",x"20",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00")



);


type object_form4 is array (0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic;
constant object4 : object_form4 := (
("00000000000000000000"),
("00000000000000000000"),
("00000000000000000000"),
("00000000000000011000"),
("00010000000000111100"),
("00011100000000111100"),
("00011110000001111100"),
("00011110000001111100"),
("00111110000001111100"),
("00111110000001111100"),
("00111110000001111100"),
("00111110000001111100"),
("00111110000001111100"),
("00111110000001111100"),
("00111111111111111100"),
("00111111111111111100"),
("00001111111111110000"),
("00000111111111111000"),
("00000000011111111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111000"),
("00000000000001111000"),
("00000000000001111000"),
("00000000000001111000"),
("00000000000001111000"),
("00000000000001111000"),
("00000000000000111000"),
("00000000000000000000"),
("00000000000000000000"),
("00000000000000000000")
);

type ram_array5 is array(0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic_vector(7 downto 0);
constant object_colors5: ram_array5 := ( 
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"64",x"a4",x"c4",x"a4",x"a4",x"a4",x"a4",x"84",x"84",x"84",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"a4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"64",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"20",x"20",x"60",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"a4",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"c8",x"c4",x"40",x"00",x"40",x"64",x"64",x"64",x"64",x"64",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"e8",x"e8",x"e8",x"a4",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"e8",x"e8",x"e8",x"c4",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"20",x"e8",x"e8",x"e8",x"a4",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"20",x"e8",x"e8",x"e8",x"a4",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"40",x"e8",x"e8",x"e8",x"84",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"40",x"e8",x"e8",x"e8",x"84",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"60",x"e8",x"e8",x"e8",x"64",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"64",x"e8",x"e8",x"e8",x"60",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"84",x"e8",x"e8",x"a4",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"40",x"a4",x"40",x"20",x"a4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"a4",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"60",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"40",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"40",x"c4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"84",x"20",x"20",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"64",x"c4",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"c4",x"e8",x"e8",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"c4",x"e8",x"e8",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"c4",x"e8",x"e8",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"c8",x"e8",x"e8",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"e8",x"e8",x"e8",x"e8",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"e8",x"e8",x"e8",x"e8",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"e8",x"e8",x"e8",x"e8",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"e8",x"e8",x"e8",x"c4",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"c4",x"e8",x"e8",x"c4",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"20",x"a4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"84",x"40",x"e8",x"e8",x"84",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"a4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"40",x"a4",x"c8",x"20",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"20",x"84",x"a4",x"a4",x"a4",x"a4",x"c4",x"c4",x"c4",x"c4",x"84",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00")


);


type object_form5 is array (0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic;
constant object5 : object_form5 := (
("00000000000000000000"),
("00000000000000000000"),
("00000111111111100000"),
("00001111111111100000"),
("00011111111111000000"),
("00011101111110000000"),
("00011110000000000000"),
("00011110000000000000"),
("00111110000000000000"),
("00111110000000000000"),
("00111110000000000000"),
("00111110000000000000"),
("00111110000000000000"),
("00111110000000000000"),
("00111111111110000000"),
("00111111111111000000"),
("00001111111111110000"),
("00000111111111111000"),
("00000000011111111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111000"),
("00000000000001111000"),
("00000000000001111000"),
("00000000000001111000"),
("00000011111101111000"),
("00001111111111111000"),
("00011111111111111000"),
("00011111111111000000"),
("00000000000000000000"),
("00000000000000000000")

);

type ram_array6 is array(0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic_vector(7 downto 0);
constant object_colors6: ram_array6 := ( 

(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"64",x"a4",x"c4",x"a4",x"a4",x"a4",x"a4",x"84",x"84",x"84",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"a4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"64",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"20",x"20",x"60",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"a4",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"c8",x"c4",x"40",x"00",x"40",x"64",x"64",x"64",x"64",x"64",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"e8",x"e8",x"e8",x"a4",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"e8",x"e8",x"e8",x"c4",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"20",x"e8",x"e8",x"e8",x"a4",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"20",x"e8",x"e8",x"e8",x"a4",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"40",x"e8",x"e8",x"e8",x"84",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"40",x"e8",x"e8",x"e8",x"84",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"60",x"e8",x"e8",x"e8",x"64",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"64",x"e8",x"e8",x"e8",x"60",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"84",x"e8",x"e8",x"a4",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"40",x"a4",x"40",x"20",x"a4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"a4",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"60",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"40",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"40",x"20",x"40",x"c4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"84",x"20",x"20",x"00",x"00",x"00"),
(x"00",x"00",x"64",x"e8",x"e8",x"64",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"64",x"c4",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"84",x"e8",x"e8",x"e8",x"40",x"00",x"00",x"00",x"00",x"00",x"00",x"c4",x"e8",x"e8",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"84",x"e8",x"e8",x"e8",x"40",x"00",x"00",x"00",x"00",x"00",x"00",x"c4",x"e8",x"e8",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"84",x"e8",x"e8",x"e8",x"40",x"00",x"00",x"00",x"00",x"00",x"00",x"c4",x"e8",x"e8",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"84",x"e8",x"e8",x"e8",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"c8",x"e8",x"e8",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"a4",x"e8",x"e8",x"e8",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"e8",x"e8",x"e8",x"e8",x"00",x"00",x"00"),
(x"00",x"00",x"a4",x"e8",x"e8",x"e8",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"e8",x"e8",x"e8",x"e8",x"00",x"00",x"00"),
(x"00",x"00",x"a4",x"e8",x"e8",x"e8",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"e8",x"e8",x"e8",x"e8",x"00",x"00",x"00"),
(x"00",x"00",x"a4",x"e8",x"e8",x"e8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"e8",x"e8",x"e8",x"c4",x"00",x"00",x"00"),
(x"00",x"00",x"a4",x"e8",x"a4",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"c4",x"e8",x"e8",x"c4",x"00",x"00",x"00"),
(x"00",x"00",x"64",x"40",x"20",x"a4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"84",x"40",x"e8",x"e8",x"84",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"84",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"40",x"a4",x"c8",x"20",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"20",x"84",x"a4",x"a4",x"a4",x"a4",x"c4",x"c4",x"c4",x"c4",x"84",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00")


);


type object_form6 is array (0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic;
constant object6 : object_form6 := (
("00000000000000000000"),
("00000000000000000000"),
("00000111111111100000"),
("00001111111111100000"),
("00011111111111000000"),
("00011101111110000000"),
("00011110000000000000"),
("00011110000000000000"),
("00111110000000000000"),
("00111110000000000000"),
("00111110000000000000"),
("00111110000000000000"),
("00111110000000000000"),
("00111110000000000000"),
("00111111111110000000"),
("00111111111111000000"),
("00001111111111110000"),
("00011111111111111000"),
("00111100011111111100"),
("00111110000001111100"),
("00111110000001111100"),
("00111110000001111100"),
("00111110000001111100"),
("00111110000001111000"),
("00111110000001111000"),
("00111110000001111000"),
("00111100000001111000"),
("00111111111101111000"),
("00111111111111111000"),
("00011111111111111000"),
("00011111111111000000"),
("00000000000000000000"),
("00000000000000000000")
);

type ram_array7 is array(0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic_vector(7 downto 0);
constant object_colors7: ram_array7 := ( 

(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"64",x"a4",x"c4",x"a4",x"a4",x"a4",x"a4",x"84",x"84",x"84",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"a4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"64",x"64",x"a4",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"64",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"a4",x"20",x"e8",x"e8",x"64",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"64",x"64",x"64",x"64",x"60",x"20",x"c4",x"e8",x"e8",x"a4",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"e8",x"e8",x"e8",x"a4",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"e8",x"e8",x"e8",x"84",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"e8",x"e8",x"e8",x"84",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"e8",x"e8",x"e8",x"84",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"60",x"e8",x"e8",x"e8",x"64",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"64",x"e8",x"e8",x"e8",x"60",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"64",x"e8",x"e8",x"e8",x"40",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"84",x"e8",x"e8",x"e8",x"40",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"c4",x"e8",x"e8",x"40",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"84",x"c4",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"84",x"c4",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"c4",x"e8",x"e8",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"c4",x"e8",x"e8",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"c4",x"e8",x"e8",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"c8",x"e8",x"e8",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"e8",x"e8",x"e8",x"e8",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"e8",x"e8",x"e8",x"e8",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"e8",x"e8",x"e8",x"e8",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"e8",x"e8",x"e8",x"c4",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"c4",x"e8",x"e8",x"c4",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"e8",x"e8",x"84",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"a4",x"c8",x"20",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00")

);


type object_form7 is array (0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic;
constant object7 : object_form7 := (
("00000000000000000000"),
("00000000000000000000"),
("00000111111111100000"),
("00001111111111111000"),
("00000111111111111100"),
("00000001111111111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000000011100"),
("00000000000000000000"),
("00000000000000001000"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111000"),
("00000000000001111000"),
("00000000000001111000"),
("00000000000001111000"),
("00000000000001111000"),
("00000000000001111000"),
("00000000000000111000"),
("00000000000000000000"),
("00000000000000000000"),
("00000000000000000000")

);

type ram_array8 is array(0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic_vector(7 downto 0);
constant object_colors8: ram_array8 := ( 
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"64",x"a4",x"c4",x"a4",x"a4",x"a4",x"a4",x"84",x"84",x"84",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"a4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"64",x"64",x"a4",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"20",x"20",x"60",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"a4",x"20",x"e8",x"e8",x"64",x"00",x"00"),
(x"00",x"00",x"00",x"c8",x"c4",x"40",x"00",x"40",x"64",x"64",x"64",x"64",x"60",x"20",x"c4",x"e8",x"e8",x"a4",x"00",x"00"),
(x"00",x"00",x"00",x"e8",x"e8",x"e8",x"a4",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"e8",x"e8",x"e8",x"a4",x"00",x"00"),
(x"00",x"00",x"00",x"e8",x"e8",x"e8",x"c4",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"e8",x"e8",x"e8",x"84",x"00",x"00"),
(x"00",x"00",x"20",x"e8",x"e8",x"e8",x"a4",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"e8",x"e8",x"e8",x"84",x"00",x"00"),
(x"00",x"00",x"20",x"e8",x"e8",x"e8",x"a4",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"e8",x"e8",x"e8",x"84",x"00",x"00"),
(x"00",x"00",x"40",x"e8",x"e8",x"e8",x"84",x"00",x"00",x"00",x"00",x"00",x"00",x"60",x"e8",x"e8",x"e8",x"64",x"00",x"00"),
(x"00",x"00",x"40",x"e8",x"e8",x"e8",x"84",x"00",x"00",x"00",x"00",x"00",x"00",x"64",x"e8",x"e8",x"e8",x"60",x"00",x"00"),
(x"00",x"00",x"60",x"e8",x"e8",x"e8",x"64",x"00",x"00",x"00",x"00",x"00",x"00",x"64",x"e8",x"e8",x"e8",x"40",x"00",x"00"),
(x"00",x"00",x"64",x"e8",x"e8",x"e8",x"60",x"00",x"00",x"00",x"00",x"00",x"00",x"84",x"e8",x"e8",x"e8",x"40",x"00",x"00"),
(x"00",x"00",x"84",x"e8",x"e8",x"a4",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"c4",x"e8",x"e8",x"40",x"00",x"00"),
(x"00",x"00",x"40",x"a4",x"40",x"20",x"a4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"84",x"20",x"64",x"c4",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"60",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"40",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"40",x"20",x"40",x"c4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"84",x"20",x"20",x"00",x"00",x"00"),
(x"00",x"00",x"64",x"e8",x"e8",x"64",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"64",x"c4",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"84",x"e8",x"e8",x"e8",x"40",x"00",x"00",x"00",x"00",x"00",x"00",x"c4",x"e8",x"e8",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"84",x"e8",x"e8",x"e8",x"40",x"00",x"00",x"00",x"00",x"00",x"00",x"c4",x"e8",x"e8",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"84",x"e8",x"e8",x"e8",x"40",x"00",x"00",x"00",x"00",x"00",x"00",x"c4",x"e8",x"e8",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"84",x"e8",x"e8",x"e8",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"c8",x"e8",x"e8",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"a4",x"e8",x"e8",x"e8",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"e8",x"e8",x"e8",x"e8",x"00",x"00",x"00"),
(x"00",x"00",x"a4",x"e8",x"e8",x"e8",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"e8",x"e8",x"e8",x"e8",x"00",x"00",x"00"),
(x"00",x"00",x"a4",x"e8",x"e8",x"e8",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"e8",x"e8",x"e8",x"e8",x"00",x"00",x"00"),
(x"00",x"00",x"a4",x"e8",x"e8",x"e8",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"e8",x"e8",x"e8",x"c4",x"00",x"00",x"00"),
(x"00",x"00",x"a4",x"e8",x"a4",x"40",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"c4",x"e8",x"e8",x"c4",x"00",x"00",x"00"),
(x"00",x"00",x"64",x"40",x"20",x"a4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"84",x"40",x"e8",x"e8",x"84",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"84",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"40",x"a4",x"c8",x"20",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"20",x"84",x"a4",x"a4",x"a4",x"a4",x"c4",x"c4",x"c4",x"c4",x"84",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00")



);


type object_form8 is array (0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic;
constant object8 : object_form8 := (
("00000000000000000000"),
("00000000000000000000"),
("00000111111111100000"),
("00001111111111111000"),
("00011111111111111100"),
("00011101111111111100"),
("00011110000001111100"),
("00011110000001111100"),
("00111110000001111100"),
("00111110000001111100"),
("00111110000001111100"),
("00111110000001111100"),
("00111110000001111100"),
("00111110000001111100"),
("00111111111111111100"),
("00111111111111111100"),
("00001111111111110000"),
("00011111111111111000"),
("00111100011111111100"),
("00111110000001111100"),
("00111110000001111100"),
("00111110000001111100"),
("00111110000001111100"),
("00111110000001111000"),
("00111110000001111000"),
("00111110000001111000"),
("00111100000001111000"),
("00111111111101111000"),
("00111111111111111000"),
("00011111111111111000"),
("00011111111111000000"),
("00000000000000000000"),
("00000000000000000000")
);

type ram_array9 is array(0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic_vector(7 downto 0);
constant object_colors9: ram_array9 := ( 

(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"64",x"a4",x"c4",x"a4",x"a4",x"a4",x"a4",x"84",x"84",x"84",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"a4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"64",x"64",x"a4",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"20",x"20",x"60",x"c8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"a4",x"20",x"e8",x"e8",x"64",x"00",x"00"),
(x"00",x"00",x"00",x"c8",x"c4",x"40",x"00",x"40",x"64",x"64",x"64",x"64",x"60",x"20",x"c4",x"e8",x"e8",x"a4",x"00",x"00"),
(x"00",x"00",x"00",x"e8",x"e8",x"e8",x"a4",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"e8",x"e8",x"e8",x"a4",x"00",x"00"),
(x"00",x"00",x"00",x"e8",x"e8",x"e8",x"c4",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"e8",x"e8",x"e8",x"84",x"00",x"00"),
(x"00",x"00",x"20",x"e8",x"e8",x"e8",x"a4",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"e8",x"e8",x"e8",x"84",x"00",x"00"),
(x"00",x"00",x"20",x"e8",x"e8",x"e8",x"a4",x"00",x"00",x"00",x"00",x"00",x"00",x"40",x"e8",x"e8",x"e8",x"84",x"00",x"00"),
(x"00",x"00",x"40",x"e8",x"e8",x"e8",x"84",x"00",x"00",x"00",x"00",x"00",x"00",x"60",x"e8",x"e8",x"e8",x"64",x"00",x"00"),
(x"00",x"00",x"40",x"e8",x"e8",x"e8",x"84",x"00",x"00",x"00",x"00",x"00",x"00",x"64",x"e8",x"e8",x"e8",x"60",x"00",x"00"),
(x"00",x"00",x"60",x"e8",x"e8",x"e8",x"64",x"00",x"00",x"00",x"00",x"00",x"00",x"64",x"e8",x"e8",x"e8",x"40",x"00",x"00"),
(x"00",x"00",x"64",x"e8",x"e8",x"e8",x"60",x"00",x"00",x"00",x"00",x"00",x"00",x"84",x"e8",x"e8",x"e8",x"40",x"00",x"00"),
(x"00",x"00",x"84",x"e8",x"e8",x"a4",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"c4",x"e8",x"e8",x"40",x"00",x"00"),
(x"00",x"00",x"40",x"a4",x"40",x"20",x"a4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"84",x"20",x"64",x"c4",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"60",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"40",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"40",x"c4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"c4",x"84",x"20",x"20",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"64",x"c4",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"c4",x"e8",x"e8",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"c4",x"e8",x"e8",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"c4",x"e8",x"e8",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"c8",x"e8",x"e8",x"e8",x"20",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"e8",x"e8",x"e8",x"e8",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"e8",x"e8",x"e8",x"e8",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"e8",x"e8",x"e8",x"e8",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"e8",x"e8",x"e8",x"c4",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"20",x"20",x"20",x"00",x"c4",x"e8",x"e8",x"c4",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"20",x"a4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"84",x"40",x"e8",x"e8",x"84",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"a4",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"e8",x"40",x"a4",x"c8",x"20",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"20",x"84",x"a4",x"a4",x"a4",x"a4",x"c4",x"c4",x"c4",x"c4",x"84",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"),
(x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00")


);


type object_form9 is array (0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic;
constant object9 : object_form9 := (
("00000000000000000000"),
("00000000000000000000"),
("00000111111111100000"),
("00001111111111111000"),
("00011111111111111100"),
("00011101111111111100"),
("00011110000001111100"),
("00011110000001111100"),
("00111110000001111100"),
("00111110000001111100"),
("00111110000001111100"),
("00111110000001111100"),
("00111110000001111100"),
("00111110000001111100"),
("00111111111111111100"),
("00111111111111111100"),
("00001111111111110000"),
("00000111111111111000"),
("00000000011111111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111100"),
("00000000000001111000"),
("00000000000001111000"),
("00000000000001111000"),
("00000000000001111000"),
("00000011111101111000"),
("00001111111111111000"),
("00011111111111111000"),
("00011111111111000000"),
("00000000000000000000"),
("00000000000000000000")
);


signal  LSB_number  : integer := 0;

signal bCoord_X : integer := 0;-- offset from start position 
signal bCoord_Y : integer := 0;

signal drawing_X : std_logic := '0';
signal drawing_Y : std_logic := '0';

--		
signal objectEndX : integer;
signal objectEndY : integer;

begin


-- Calculate object end boundaries
objectEndX	<= object_X_size+ObjectStartX;
objectEndY	<= object_Y_size+ObjectStartY;


-- Signals drawing_X[Y] are active when obects coordinates are being crossed

-- test if ooCoord is in the rectangle defined by Start and End 
	drawing_X	<= '1' when  (oCoord_X  >= ObjectStartX) and  (oCoord_X < objectEndX) else '0';
    drawing_Y	<= '1' when  (oCoord_Y  >= ObjectStartY) and  (oCoord_Y < objectEndY) else '0';
	 

	bCoord_X 	<= (oCoord_X - ObjectStartX) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 
	bCoord_Y 	<= (oCoord_Y - ObjectStartY) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 


process ( RESETn, CLK)

   begin
	
	if RESETn = '0' then
	    mVGA_RGB	<=  (others => '0') ; 	
		drawing_request	<=  '0' ;
	     
		elsif rising_edge(CLK) then
		   
                
		      case LSB_number is 
				  when 0 => 
				    mVGA_RGB	<=  object_colors0(bCoord_Y , bCoord_X);	--get from colors table 
			       drawing_request	<= object0(bCoord_Y , bCoord_X) and drawing_X and drawing_Y ; -- get from mask table 	
				  when 1 => 
				    mVGA_RGB	<=  object_colors1(bCoord_Y , bCoord_X);	--get from colors table 
			       drawing_request	<= object1(bCoord_Y , bCoord_X) and drawing_X and drawing_Y ; -- get from mask table 	 	
 				  when 2 => 
				    mVGA_RGB	<=  object_colors2(bCoord_Y , bCoord_X);	--get from colors table 
			       drawing_request	<= object2(bCoord_Y , bCoord_X) and drawing_X and drawing_Y ; -- get from mask table 
				  when 3 => 
				    mVGA_RGB	<=  object_colors3(bCoord_Y , bCoord_X);	--get from colors table 
			       drawing_request	<= object3(bCoord_Y , bCoord_X) and drawing_X and drawing_Y ; -- get from mask table 	
				  when 4 => 
				    mVGA_RGB	<=  object_colors4(bCoord_Y , bCoord_X);	--get from colors table 
			       drawing_request	<= object4(bCoord_Y , bCoord_X) and drawing_X and drawing_Y ; -- get from mask table 	 
				  when 5 => 
				    mVGA_RGB	<=  object_colors5(bCoord_Y , bCoord_X);	--get from colors table 
			       drawing_request	<= object5(bCoord_Y , bCoord_X) and drawing_X and drawing_Y ; -- get from mask table 	
				  when 6 => 
				    mVGA_RGB	<=  object_colors6(bCoord_Y , bCoord_X);	--get from colors table 
			       drawing_request	<= object6(bCoord_Y , bCoord_X) and drawing_X and drawing_Y ; -- get from mask table 	
				  when 7 => 
				    mVGA_RGB	<=  object_colors7(bCoord_Y , bCoord_X);	--get from colors table 
			       drawing_request	<= object7(bCoord_Y , bCoord_X) and drawing_X and drawing_Y ; -- get from mask table 	
				  when 8 => 
				    mVGA_RGB	<=  object_colors8(bCoord_Y , bCoord_X);	--get from colors table 
			       drawing_request	<= object8(bCoord_Y , bCoord_X) and drawing_X and drawing_Y ; -- get from mask table 	
				  when 9 => 
				    mVGA_RGB	<=  object_colors9(bCoord_Y , bCoord_X);	--get from colors table 
			       drawing_request	<= object9(bCoord_Y , bCoord_X) and drawing_X and drawing_Y ; -- get from mask table 	 
               when others => drawing_request <= '0' ;
				  end case ;
					
				  			  
	 end if;
	  	

  end process;

		
end behav;		
		