--------------------------------------
-- SinTable.vhd
-- Written by Gadi and Eran Tuchman.
-- All rights reserved, Copyright 2009
--------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all ;

entity Explosion_Sound2 is
port(
  CLK     					: in std_logic;
  resetN 					: in std_logic;
  ENA                   : in std_logic;
  ADDR    					: in std_logic_vector(14 downto 0);
  Q       					: out std_logic_vector(15 downto 0)
);
end Explosion_Sound2;

architecture arch of Explosion_Sound2 is
constant array_size 			: integer := 21381 ;

type table_type is array(0 to array_size - 1) of std_logic_vector(15 downto 0);
signal sin_table				: table_type;
signal Q_tmp       			:  std_logic_vector(15 downto 0) ;



begin
 
   
  sintable_proc: process(resetN, CLK)
    constant sin_table : table_type := (
---start 0 v

X"007D",
X"0000",
X"0000",
X"007D",
X"0000",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"007D",
X"0000",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"FE89",
X"FE89",
X"FE89",
X"FE0C",
X"FE89",
X"FF83",
X"FF06",
X"FE0C",
X"FF06",
X"FE0C",
X"FD8F",
X"FE0C",
X"FF83",
X"FE0C",
X"FF06",
X"00FA",
X"FE89",
X"FF06",
X"0177",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"FE89",
X"FE89",
X"FF06",
X"FD8F",
X"FF06",
X"FD12",
X"FE89",
X"0000",
X"FF06",
X"FE0C",
X"FE0C",
X"FF06",
X"FE89",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"00FA",
X"0000",
X"007D",
X"01F4",
X"0271",
X"0271",
X"0177",
X"01F4",
X"03E8",
X"007D",
X"0177",
X"02EE",
X"0177",
X"00FA",
X"01F4",
X"03E8",
X"007D",
X"02EE",
X"00FA",
X"007D",
X"00FA",
X"0000",
X"0000",
X"0000",
X"FF06",
X"007D",
X"0000",
X"FD12",
X"007D",
X"0271",
X"00FA",
X"0177",
X"01F4",
X"02EE",
X"00FA",
X"0177",
X"0465",
X"0000",
X"0271",
X"01F4",
X"0000",
X"01F4",
X"0000",
X"0271",
X"02EE",
X"02EE",
X"007D",
X"0271",
X"FF83",
X"007D",
X"0271",
X"00FA",
X"FF83",
X"007D",
X"FF06",
X"007D",
X"0000",
X"0177",
X"0271",
X"007D",
X"0271",
X"0271",
X"02EE",
X"0271",
X"036B",
X"01F4",
X"00FA",
X"0177",
X"FF83",
X"FF06",
X"FF83",
X"FF06",
X"FC95",
X"FD12",
X"FE89",
X"FD8F",
X"FC18",
X"FC95",
X"FD12",
X"FD8F",
X"FD12",
X"FF83",
X"00FA",
X"0000",
X"00FA",
X"FD8F",
X"FC95",
X"036B",
X"0000",
X"00FA",
X"0000",
X"FF83",
X"0177",
X"0177",
X"0177",
X"FB1E",
X"FF06",
X"0177",
X"FF06",
X"0271",
X"0753",
X"0000",
X"0271",
X"03E8",
X"036B",
X"04E2",
X"00FA",
X"04E2",
X"02EE",
X"02EE",
X"036B",
X"01F4",
X"FE89",
X"FC18",
X"F9A7",
X"FA24",
X"F9A7",
X"F830",
X"F92A",
X"F92A",
X"FAA1",
X"FB9B",
X"F9A7",
X"FAA1",
X"FB9B",
X"F9A7",
X"FB1E",
X"FA24",
X"FD8F",
X"FE89",
X"FC18",
X"F8AD",
X"F9A7",
X"FD12",
X"00FA",
X"FD12",
X"FC95",
X"FE89",
X"FD12",
X"00FA",
X"0177",
X"02EE",
X"03E8",
X"03E8",
X"03E8",
X"0271",
X"01F4",
X"FF06",
X"007D",
X"01F4",
X"01F4",
X"007D",
X"02EE",
X"0271",
X"02EE",
X"036B",
X"02EE",
X"03E8",
X"01F4",
X"036B",
X"036B",
X"0465",
X"036B",
X"03E8",
X"036B",
X"03E8",
X"0271",
X"0465",
X"0271",
X"03E8",
X"03E8",
X"FE89",
X"0000",
X"FF83",
X"00FA",
X"FE89",
X"FD12",
X"FD8F",
X"FE89",
X"FD8F",
X"FF06",
X"FF06",
X"FE0C",
X"FE89",
X"FD8F",
X"FE89",
X"FC95",
X"FD12",
X"FF06",
X"0000",
X"FD12",
X"FD8F",
X"FC95",
X"FB1E",
X"FAA1",
X"F9A7",
X"FB1E",
X"F9A7",
X"FAA1",
X"FE89",
X"FD12",
X"FF06",
X"FF83",
X"0000",
X"00FA",
X"FF06",
X"00FA",
X"FF06",
X"0000",
X"007D",
X"0000",
X"036B",
X"0271",
X"0465",
X"05DC",
X"0659",
X"05DC",
X"0659",
X"084D",
X"08CA",
X"055F",
X"055F",
X"055F",
X"0465",
X"02EE",
X"03E8",
X"0000",
X"0177",
X"00FA",
X"FD12",
X"FB9B",
X"FD12",
X"F92A",
X"FC95",
X"00FA",
X"FF06",
X"01F4",
X"04E2",
X"01F4",
X"007D",
X"0271",
X"01F4",
X"02EE",
X"FD8F",
X"FC18",
X"FE89",
X"FC18",
X"FD8F",
X"FC95",
X"FD8F",
X"FD8F",
X"FD8F",
X"0271",
X"FF83",
X"0000",
X"01F4",
X"FB1E",
X"FB1E",
X"FD8F",
X"0465",
X"FC18",
X"0000",
X"FF06",
X"007D",
X"FF83",
X"FB1E",
X"FF06",
X"FD12",
X"FF06",
X"FE0C",
X"FF83",
X"FE89",
X"FE89",
X"00FA",
X"FC18",
X"FE0C",
X"FC18",
X"FF83",
X"FE0C",
X"FA24",
X"F5BF",
X"FAA1",
X"F63C",
X"F9A7",
X"F9A7",
X"F448",
X"FA24",
X"FB9B",
X"FD12",
X"F7B3",
X"FE89",
X"0000",
X"FD12",
X"0000",
X"06D6",
X"FAA1",
X"0947",
X"0FA0",
X"05DC",
X"16F3",
X"0B3B",
X"130B",
X"16F3",
X"109A",
X"0E29",
X"0BB8",
X"0ABE",
X"0947",
X"09C4",
X"128E",
X"FE89",
X"1117",
X"0177",
X"0D2F",
X"0659",
X"EA07",
X"FD8F",
X"F5BF",
X"F4C5",
X"F3CB",
X"FC18",
X"07D0",
X"F7B3",
X"1B58",
X"0000",
X"007D",
X"F8AD",
X"08CA",
X"18E7",
X"128E",
X"1EC3",
X"09C4",
X"084D",
X"06D6",
X"F2D1",
X"03E8",
X"E98A",
X"FC95",
X"ECF5",
X"ECF5",
X"F6B9",
X"E813",
X"DC5B",
X"E90D",
X"E813",
X"E42B",
X"E1BA",
X"E719",
X"F060",
X"FAA1",
X"FB9B",
X"1388",
X"09C4",
X"F254",
X"F3CB",
X"0947",
X"007D",
X"F34E",
X"F3CB",
X"0271",
X"1770",
X"130B",
X"1194",
X"0659",
X"06D6",
X"0CB2",
X"1117",
X"0947",
X"09C4",
X"036B",
X"02EE",
X"F2D1",
X"F4C5",
X"FC95",
X"EBFB",
X"EEE9",
X"EE6C",
X"EA84",
X"E5A2",
X"E043",
X"D873",
X"CA4A",
X"C662",
X"CA4A",
X"CBC1",
X"D19D",
X"D7F6",
X"ECF5",
X"F5BF",
X"E3AE",
X"FD8F",
X"130B",
X"09C4",
X"04E2",
X"2422",
X"1C52",
X"1ADB",
X"20B7",
X"1D4C",
X"203A",
X"1D4C",
X"0E29",
X"101D",
X"1FBD",
X"FAA1",
X"0947",
X"1211",
X"F9A7",
X"0659",
X"ECF5",
X"07D0",
X"0753",
X"06D6",
X"FE0C",
X"F1D7",
X"FAA1",
X"F63C",
X"FB9B",
X"06D6",
X"FD12",
X"09C4",
X"203A",
X"0ABE",
X"1117",
X"1ADB",
X"1E46",
X"2B75",
X"3539",
X"31CE",
X"251C",
X"22AB",
X"37AA",
X"3151",
X"2A7B",
X"2599",
X"20B7",
X"0EA6",
X"0659",
X"1ADB",
X"18E7",
X"0CB2",
X"0B3B",
X"0753",
X"F15A",
X"FD8F",
X"0C35",
X"0000",
X"FA24",
X"ECF5",
X"F448",
X"DFC6",
X"E90D",
X"EC78",
X"EC78",
X"F2D1",
X"F5BF",
X"05DC",
X"1211",
X"1676",
X"17ED",
X"18E7",
X"1405",
X"1211",
X"1117",
X"09C4",
X"0177",
X"EEE9",
X"F830",
X"FD12",
X"F34E",
X"F542",
X"EE6C",
X"ECF5",
X"E98A",
X"E69C",
X"E69C",
X"E42B",
X"E525",
X"E61F",
X"E4A8",
X"E61F",
X"E796",
X"E13D",
X"CF2C",
X"D0A3",
X"D67F",
X"D67F",
X"EE6C",
X"F254",
X"F0DD",
X"F3CB",
X"F830",
X"F830",
X"F830",
X"F2D1",
X"E2B4",
X"F34E",
X"F9A7",
X"F63C",
X"F830",
X"F92A",
X"FA24",
X"F736",
X"F542",
X"F830",
X"F736",
X"F448",
X"F6B9",
X"F0DD",
X"F34E",
X"F63C",
X"FB1E",
X"FC95",
X"FB9B",
X"FB1E",
X"F7B3",
X"F542",
X"EA07",
X"EEE9",
X"EFE3",
X"F63C",
X"F830",
X"F542",
X"02EE",
X"07D0",
X"0F23",
X"14FF",
X"130B",
X"1676",
X"1D4C",
X"1EC3",
X"21B1",
X"2616",
X"20B7",
X"2616",
X"2328",
X"2BF2",
X"2E63",
X"1FBD",
X"2981",
X"1BD5",
X"1D4C",
X"1C52",
X"16F3",
X"1676",
X"1117",
X"109A",
X"0BB8",
X"0465",
X"08CA",
X"03E8",
X"02EE",
X"FC18",
X"FD12",
X"F830",
X"F63C",
X"F92A",
X"F254",
X"F15A",
X"F060",
X"F4C5",
X"F254",
X"FC18",
X"F8AD",
X"FF83",
X"055F",
X"FF06",
X"0177",
X"01F4",
X"007D",
X"FAA1",
X"FB9B",
X"F736",
X"F3CB",
X"E90D",
X"E890",
X"DE4F",
X"D297",
X"DA67",
X"E719",
X"DAE4",
X"D67F",
X"DB61",
X"D6FC",
X"E3AE",
X"E2B4",
X"ECF5",
X"E61F",
X"E2B4",
X"FC95",
X"F830",
X"01F4",
X"FD12",
X"FB9B",
X"0271",
X"05DC",
X"00FA",
X"036B",
X"055F",
X"FE89",
X"007D",
X"FF06",
X"FC95",
X"FC95",
X"F9A7",
X"FE89",
X"01F4",
X"0271",
X"0271",
X"00FA",
X"0271",
X"09C4",
X"06D6",
X"02EE",
X"07D0",
X"0CB2",
X"084D",
X"07D0",
X"09C4",
X"0A41",
X"0EA6",
X"0EA6",
X"128E",
X"109A",
X"130B",
X"1388",
X"0DAC",
X"19E1",
X"1482",
X"0F23",
X"1482",
X"15F9",
X"0EA6",
X"06D6",
X"0B3B",
X"1482",
X"109A",
X"14FF",
X"128E",
X"1211",
X"186A",
X"20B7",
X"1FBD",
X"2693",
X"22AB",
X"2887",
X"2599",
X"2A7B",
X"251C",
X"2887",
X"2887",
X"20B7",
X"2710",
X"22AB",
X"2134",
X"2616",
X"22AB",
X"22AB",
X"2328",
X"1ADB",
X"16F3",
X"128E",
X"14FF",
X"1117",
X"0947",
X"0B3B",
X"07D0",
X"0753",
X"0BB8",
X"FF06",
X"01F4",
X"0465",
X"03E8",
X"FE89",
X"F2D1",
X"F736",
X"ED72",
X"E890",
X"E2B4",
X"DFC6",
X"E13D",
X"E237",
X"E796",
X"EDEF",
X"EB7E",
X"F0DD",
X"E813",
X"E90D",
X"EA84",
X"E719",
X"E61F",
X"E13D",
X"E69C",
X"E237",
X"DD55",
X"DB61",
X"DDD2",
X"DA67",
X"D585",
X"D7F6",
X"DB61",
X"D508",
X"D21A",
X"D7F6",
X"D120",
X"CC3E",
X"CBC1",
X"CA4A",
X"CC3E",
X"CF2C",
X"D96D",
X"D6FC",
X"E525",
X"EC78",
X"E1BA",
X"E237",
X"E796",
X"F15A",
X"EDEF",
X"F060",
X"FC95",
X"FF06",
X"01F4",
X"05DC",
X"109A",
X"16F3",
X"203A",
X"2CEC",
X"3345",
X"32C8",
X"2E63",
X"3057",
X"2CEC",
X"249F",
X"22AB",
X"1964",
X"1211",
X"0271",
X"F3CB",
X"FE89",
X"F254",
X"EB7E",
X"EEE9",
X"ED72",
X"FB1E",
X"FA24",
X"F9A7",
X"F060",
X"EE6C",
X"EFE3",
X"EF66",
X"F2D1",
X"F4C5",
X"F830",
X"FC95",
X"0C35",
X"109A",
X"128E",
X"14FF",
X"1405",
X"0E29",
X"09C4",
X"07D0",
X"036B",
X"06D6",
X"06D6",
X"0C35",
X"06D6",
X"036B",
X"0B3B",
X"05DC",
X"07D0",
X"101D",
X"1ADB",
X"2134",
X"1F40",
X"1EC3",
X"222E",
X"1FBD",
X"1CCF",
X"128E",
X"1211",
X"0FA0",
X"09C4",
X"0947",
X"0000",
X"FAA1",
X"F448",
X"F5BF",
X"EFE3",
X"E69C",
X"E1BA",
X"DECC",
X"DD55",
X"E0C0",
X"E331",
X"E98A",
X"F448",
X"F92A",
X"F5BF",
X"F8AD",
X"EF66",
X"F0DD",
X"EF66",
X"EA07",
X"F4C5",
X"FA24",
X"01F4",
X"0271",
X"FC18",
X"01F4",
X"0465",
X"03E8",
X"08CA",
X"0E29",
X"1BD5",
X"1A5E",
X"1194",
X"0947",
X"1405",
X"1770",
X"2134",
X"2710",
X"249F",
X"2C6F",
X"30D4",
X"1FBD",
X"17ED",
X"109A",
X"1211",
X"0ABE",
X"084D",
X"05DC",
X"FE89",
X"0465",
X"FF06",
X"FD8F",
X"FC95",
X"FAA1",
X"F2D1",
X"FC95",
X"F5BF",
X"FC18",
X"FB1E",
X"F4C5",
X"F7B3",
X"F254",
X"F448",
X"EF66",
X"EDEF",
X"F5BF",
X"0177",
X"FE89",
X"F5BF",
X"EE6C",
X"F15A",
X"EC78",
X"E90D",
X"EBFB",
X"E890",
X"E890",
X"EFE3",
X"F0DD",
X"F15A",
X"F830",
X"F6B9",
X"F63C",
X"F2D1",
X"F4C5",
X"F542",
X"F448",
X"F8AD",
X"F4C5",
X"F736",
X"F7B3",
X"F63C",
X"F92A",
X"FAA1",
X"FE0C",
X"FF06",
X"FF06",
X"FF06",
X"FAA1",
X"F92A",
X"F92A",
X"FAA1",
X"F830",
X"FB1E",
X"F736",
X"F92A",
X"FB1E",
X"FC95",
X"FB9B",
X"FB9B",
X"036B",
X"FD8F",
X"FF06",
X"FD8F",
X"FE0C",
X"F9A7",
X"FC18",
X"F8AD",
X"FD8F",
X"FE89",
X"FF06",
X"FF83",
X"01F4",
X"0C35",
X"084D",
X"0E29",
X"109A",
X"109A",
X"1211",
X"130B",
X"109A",
X"101D",
X"1388",
X"0BB8",
X"0CB2",
X"0A41",
X"0D2F",
X"0E29",
X"0DAC",
X"1117",
X"084D",
X"09C4",
X"0CB2",
X"01F4",
X"0D2F",
X"0465",
X"0659",
X"0A41",
X"07D0",
X"06D6",
X"0659",
X"036B",
X"0659",
X"08CA",
X"0000",
X"FF06",
X"0659",
X"FB1E",
X"FF06",
X"0000",
X"F4C5",
X"F542",
X"F2D1",
X"F3CB",
X"EA07",
X"EBFB",
X"EC78",
X"EC78",
X"EEE9",
X"EBFB",
X"EB01",
X"F542",
X"F2D1",
X"FD8F",
X"F92A",
X"FA24",
X"FB1E",
X"FD8F",
X"FF06",
X"F7B3",
X"F9A7",
X"FE89",
X"F5BF",
X"FF06",
X"FB9B",
X"FC95",
X"007D",
X"FE0C",
X"02EE",
X"0177",
X"FE89",
X"FB9B",
X"FF06",
X"FB9B",
X"03E8",
X"00FA",
X"0177",
X"00FA",
X"FE0C",
X"0000",
X"FD8F",
X"FF06",
X"0465",
X"0D2F",
X"0BB8",
X"0B3B",
X"1405",
X"0A41",
X"1388",
X"109A",
X"0FA0",
X"1194",
X"109A",
X"1194",
X"0E29",
X"0E29",
X"0FA0",
X"101D",
X"101D",
X"0C35",
X"0DAC",
X"0D2F",
X"0C35",
X"0ABE",
X"0DAC",
X"0CB2",
X"0947",
X"0BB8",
X"0753",
X"0A41",
X"055F",
X"0BB8",
X"0659",
X"0ABE",
X"0D2F",
X"0659",
X"0B3B",
X"07D0",
X"1194",
X"0DAC",
X"0E29",
X"1388",
X"1211",
X"0E29",
X"0FA0",
X"1388",
X"109A",
X"109A",
X"0BB8",
X"128E",
X"0F23",
X"0DAC",
X"0F23",
X"0B3B",
X"09C4",
X"0465",
X"06D6",
X"0465",
X"0177",
X"FF83",
X"FF06",
X"F8AD",
X"FE89",
X"FB9B",
X"FB1E",
X"FE89",
X"F8AD",
X"FD8F",
X"FA24",
X"FD12",
X"FE89",
X"FE0C",
X"FF06",
X"FAA1",
X"FC18",
X"FC18",
X"F8AD",
X"FA24",
X"F736",
X"F3CB",
X"EF66",
X"F060",
X"E90D",
X"E796",
X"E719",
X"E719",
X"E525",
X"E3AE",
X"E1BA",
X"E61F",
X"E796",
X"E796",
X"EB7E",
X"E90D",
X"EA84",
X"EF66",
X"EB01",
X"EE6C",
X"EFE3",
X"EE6C",
X"F254",
X"F2D1",
X"F5BF",
X"F7B3",
X"FA24",
X"F830",
X"F448",
X"F4C5",
X"F7B3",
X"F34E",
X"F15A",
X"F736",
X"F7B3",
X"F736",
X"F92A",
X"F542",
X"F8AD",
X"F542",
X"F9A7",
X"F5BF",
X"FA24",
X"FB1E",
X"FA24",
X"01F4",
X"007D",
X"0465",
X"0465",
X"04E2",
X"08CA",
X"0659",
X"0947",
X"055F",
X"0753",
X"04E2",
X"0947",
X"02EE",
X"0000",
X"00FA",
X"FF06",
X"0177",
X"FF83",
X"01F4",
X"03E8",
X"03E8",
X"00FA",
X"FD8F",
X"FC18",
X"FF06",
X"F830",
X"FC95",
X"F736",
X"F7B3",
X"F6B9",
X"FF83",
X"FB9B",
X"EA07",
X"EE6C",
X"ECF5",
X"F2D1",
X"FAA1",
X"EB7E",
X"F736",
X"F15A",
X"EC78",
X"F060",
X"EE6C",
X"EEE9",
X"EEE9",
X"F5BF",
X"F63C",
X"F7B3",
X"F9A7",
X"FF83",
X"0271",
X"007D",
X"0271",
X"055F",
X"055F",
X"0B3B",
X"0947",
X"0B3B",
X"0FA0",
X"0F23",
X"15F9",
X"1211",
X"128E",
X"15F9",
X"16F3",
X"186A",
X"19E1",
X"14FF",
X"130B",
X"1B58",
X"18E7",
X"278D",
X"1EC3",
X"14FF",
X"1676",
X"1117",
X"0E29",
X"0D2F",
X"109A",
X"08CA",
X"0B3B",
X"0659",
X"0659",
X"01F4",
X"07D0",
X"0271",
X"00FA",
X"FE0C",
X"007D",
X"FF06",
X"FD8F",
X"00FA",
X"F63C",
X"FAA1",
X"FC18",
X"FB1E",
X"F4C5",
X"FD8F",
X"0271",
X"FD12",
X"084D",
X"00FA",
X"0659",
X"05DC",
X"F9A7",
X"0B3B",
X"02EE",
X"0BB8",
X"05DC",
X"007D",
X"0465",
X"0177",
X"07D0",
X"0947",
X"0A41",
X"055F",
X"0465",
X"01F4",
X"FE0C",
X"FD12",
X"F1D7",
X"F63C",
X"F4C5",
X"F1D7",
X"F254",
X"EDEF",
X"E796",
X"F1D7",
X"ED72",
X"EC78",
X"EE6C",
X"EBFB",
X"EFE3",
X"F1D7",
X"F2D1",
X"F7B3",
X"F2D1",
X"F8AD",
X"0BB8",
X"FB1E",
X"F830",
X"0A41",
X"FB9B",
X"0753",
X"01F4",
X"FC95",
X"007D",
X"F92A",
X"0D2F",
X"07D0",
X"FB1E",
X"055F",
X"06D6",
X"055F",
X"F6B9",
X"FE0C",
X"F9A7",
X"F63C",
X"F254",
X"FF06",
X"036B",
X"FC18",
X"0ABE",
X"09C4",
X"FC18",
X"FF06",
X"FB9B",
X"FD8F",
X"F4C5",
X"F92A",
X"F830",
X"F254",
X"F4C5",
X"F7B3",
X"FD12",
X"F542",
X"07D0",
X"0C35",
X"0000",
X"0465",
X"F5BF",
X"0753",
X"06D6",
X"0ABE",
X"0947",
X"036B",
X"09C4",
X"0B3B",
X"0B3B",
X"0753",
X"0947",
X"0CB2",
X"0CB2",
X"0947",
X"0A41",
X"0CB2",
X"00FA",
X"05DC",
X"036B",
X"FC95",
X"055F",
X"0465",
X"00FA",
X"FF83",
X"01F4",
X"FC18",
X"00FA",
X"FC95",
X"FE0C",
X"0177",
X"055F",
X"0947",
X"FE89",
X"F5BF",
X"F542",
X"FC18",
X"FB1E",
X"FF83",
X"FB9B",
X"036B",
X"07D0",
X"0465",
X"15F9",
X"0CB2",
X"130B",
X"1194",
X"0A41",
X"14FF",
X"101D",
X"101D",
X"1117",
X"0ABE",
X"0EA6",
X"0DAC",
X"036B",
X"08CA",
X"04E2",
X"007D",
X"0659",
X"FD12",
X"007D",
X"007D",
X"FB9B",
X"FD12",
X"F63C",
X"F7B3",
X"F3CB",
X"F34E",
X"EEE9",
X"F15A",
X"F92A",
X"F2D1",
X"F15A",
X"ED72",
X"FAA1",
X"F9A7",
X"EB01",
X"F2D1",
X"00FA",
X"E4A8",
X"EEE9",
X"F34E",
X"F060",
X"FF83",
X"FD12",
X"109A",
X"05DC",
X"FF06",
X"0CB2",
X"08CA",
X"0FA0",
X"0D2F",
X"0F23",
X"1117",
X"128E",
X"1ADB",
X"20B7",
X"1A5E",
X"0BB8",
X"0CB2",
X"0FA0",
X"084D",
X"06D6",
X"0DAC",
X"0659",
X"0F23",
X"0B3B",
X"09C4",
X"1964",
X"007D",
X"01F4",
X"0B3B",
X"007D",
X"055F",
X"0A41",
X"07D0",
X"0177",
X"0ABE",
X"0271",
X"00FA",
X"F4C5",
X"FD8F",
X"FB9B",
X"F8AD",
X"FD12",
X"F63C",
X"FF83",
X"F736",
X"F63C",
X"F8AD",
X"F0DD",
X"F254",
X"F2D1",
X"EF66",
X"F448",
X"F34E",
X"F1D7",
X"F9A7",
X"FA24",
X"F060",
X"F3CB",
X"F2D1",
X"FF83",
X"F34E",
X"0177",
X"07D0",
X"007D",
X"0753",
X"055F",
X"0177",
X"FD8F",
X"01F4",
X"FE0C",
X"0177",
X"FF83",
X"08CA",
X"036B",
X"06D6",
X"FF83",
X"06D6",
X"0A41",
X"0D2F",
X"084D",
X"FC18",
X"0ABE",
X"FE0C",
X"F92A",
X"FAA1",
X"F7B3",
X"F060",
X"F7B3",
X"F830",
X"0000",
X"FB1E",
X"F6B9",
X"05DC",
X"EDEF",
X"EF66",
X"F736",
X"EA07",
X"DA67",
X"E90D",
X"EBFB",
X"DCD8",
X"DC5B",
X"E043",
X"E0C0",
X"E42B",
X"E2B4",
X"E813",
X"EC78",
X"EBFB",
X"ED72",
X"ECF5",
X"ED72",
X"ECF5",
X"F3CB",
X"F3CB",
X"F060",
X"F7B3",
X"F1D7",
X"FE89",
X"0177",
X"EC78",
X"FF06",
X"FF06",
X"0177",
X"04E2",
X"F9A7",
X"0A41",
X"0B3B",
X"0A41",
X"0947",
X"01F4",
X"0FA0",
X"0BB8",
X"0DAC",
X"0E29",
X"109A",
X"1770",
X"0ABE",
X"1482",
X"1770",
X"0B3B",
X"0CB2",
X"0ABE",
X"0BB8",
X"16F3",
X"14FF",
X"20B7",
X"101D",
X"29FE",
X"20B7",
X"1CCF",
X"203A",
X"1ADB",
X"2134",
X"1D4C",
X"2C6F",
X"157C",
X"280A",
X"1EC3",
X"2328",
X"2616",
X"203A",
X"2D69",
X"22AB",
X"16F3",
X"23A5",
X"22AB",
X"1EC3",
X"109A",
X"0E29",
X"0E29",
X"02EE",
X"F8AD",
X"0659",
X"FD12",
X"0271",
X"F542",
X"FC18",
X"F1D7",
X"EDEF",
X"F254",
X"EDEF",
X"F15A",
X"ECF5",
X"E98A",
X"EBFB",
X"E90D",
X"EB7E",
X"F060",
X"F1D7",
X"EB01",
X"E42B",
X"E3AE",
X"DA67",
X"E42B",
X"E1BA",
X"F060",
X"E42B",
X"DA67",
X"DF49",
X"E13D",
X"D9EA",
X"E3AE",
X"E13D",
X"DDD2",
X"E3AE",
X"D8F0",
X"DD55",
X"D314",
X"E525",
X"D314",
X"DB61",
X"DB61",
X"E13D",
X"E719",
X"D873",
X"EA07",
X"E796",
X"DECC",
X"EF66",
X"E42B",
X"F3CB",
X"EBFB",
X"EC78",
X"E813",
X"E813",
X"ED72",
X"D67F",
X"E237",
X"E69C",
X"E3AE",
X"E813",
X"EA84",
X"EB7E",
X"F2D1",
X"EFE3",
X"F5BF",
X"FC95",
X"FAA1",
X"FD8F",
X"0F23",
X"128E",
X"0CB2",
X"0BB8",
X"0F23",
X"16F3",
X"15F9",
X"1117",
X"19E1",
X"1F40",
X"2B75",
X"2887",
X"2328",
X"2981",
X"2904",
X"29FE",
X"2C6F",
X"2F5D",
X"1CCF",
X"2904",
X"2EE0",
X"2DE6",
X"2AF8",
X"2BF2",
X"3633",
X"2E63",
X"2BF2",
X"2AF8",
X"2710",
X"2981",
X"3345",
X"3057",
X"29FE",
X"2134",
X"280A",
X"2904",
X"1964",
X"0E29",
X"1211",
X"130B",
X"F830",
X"F92A",
X"FE0C",
X"DDD2",
X"F6B9",
X"E813",
X"CF2C",
X"DC5B",
X"D19D",
X"DECC",
X"D6FC",
X"D297",
X"DCD8",
X"D8F0",
X"DC5B",
X"E90D",
X"DFC6",
X"E90D",
X"F448",
X"FB9B",
X"0000",
X"F92A",
X"F1D7",
X"F63C",
X"036B",
X"1405",
X"0C35",
X"08CA",
X"109A",
X"0EA6",
X"101D",
X"109A",
X"1211",
X"036B",
X"055F",
X"036B",
X"0177",
X"FB1E",
X"0947",
X"157C",
X"0465",
X"0271",
X"01F4",
X"FC18",
X"F6B9",
X"F2D1",
X"FB1E",
X"F7B3",
X"FE89",
X"0F23",
X"FB1E",
X"101D",
X"1405",
X"128E",
X"20B7",
X"20B7",
X"1DC9",
X"1DC9",
X"20B7",
X"2FDA",
X"2328",
X"1BD5",
X"1B58",
X"1C52",
X"128E",
X"1770",
X"0B3B",
X"101D",
X"FE89",
X"1211",
X"0BB8",
X"FE89",
X"0753",
X"01F4",
X"0947",
X"01F4",
X"01F4",
X"03E8",
X"01F4",
X"0271",
X"FF06",
X"036B",
X"0000",
X"0000",
X"F0DD",
X"0271",
X"F4C5",
X"F34E",
X"F736",
X"F0DD",
X"F9A7",
X"E98A",
X"F63C",
X"F4C5",
X"F6B9",
X"F830",
X"F448",
X"F736",
X"F830",
X"F5BF",
X"FC95",
X"FB9B",
X"F8AD",
X"F1D7",
X"F254",
X"EE6C",
X"EFE3",
X"EEE9",
X"EDEF",
X"F542",
X"EBFB",
X"0177",
X"F34E",
X"F7B3",
X"F5BF",
X"03E8",
X"084D",
X"00FA",
X"FF06",
X"FC18",
X"00FA",
X"F830",
X"06D6",
X"F63C",
X"0ABE",
X"0D2F",
X"18E7",
X"157C",
X"0465",
X"0EA6",
X"1E46",
X"1BD5",
X"0E29",
X"1BD5",
X"0ABE",
X"157C",
X"05DC",
X"0947",
X"055F",
X"FD12",
X"F1D7",
X"E1BA",
X"F060",
X"ECF5",
X"EA84",
X"DB61",
X"D40E",
X"E237",
X"E69C",
X"DAE4",
X"DFC6",
X"E043",
X"E796",
X"EC78",
X"EA84",
X"F3CB",
X"ED72",
X"EF66",
X"FC95",
X"FF83",
X"0177",
X"0C35",
X"1770",
X"18E7",
X"0947",
X"14FF",
X"1A5E",
X"1770",
X"09C4",
X"05DC",
X"0465",
X"0CB2",
X"0177",
X"FF83",
X"130B",
X"0EA6",
X"0947",
X"0C35",
X"F9A7",
X"0947",
X"F736",
X"ED72",
X"F63C",
X"ED72",
X"F542",
X"E5A2",
X"E813",
X"E4A8",
X"ECF5",
X"DC5B",
X"D9EA",
X"E890",
X"D873",
X"DBDE",
X"DFC6",
X"ECF5",
X"D9EA",
X"E796",
X"EA84",
X"E3AE",
X"F63C",
X"E525",
X"FE89",
X"E98A",
X"EE6C",
X"F1D7",
X"ED72",
X"DE4F",
X"EB01",
X"F254",
X"E890",
X"0753",
X"EF66",
X"0659",
X"0659",
X"0D2F",
X"15F9",
X"1388",
X"1964",
X"1E46",
X"1482",
X"23A5",
X"2887",
X"1D4C",
X"280A",
X"1FBD",
X"32C8",
X"2904",
X"2328",
X"2F5D",
X"2904",
X"1FBD",
X"2887",
X"2599",
X"1DC9",
X"203A",
X"1A5E",
X"1B58",
X"1E46",
X"1676",
X"15F9",
X"0FA0",
X"1964",
X"18E7",
X"0A41",
X"0EA6",
X"0000",
X"FD12",
X"FE0C",
X"F7B3",
X"F34E",
X"EB7E",
X"E237",
X"E5A2",
X"DB61",
X"DF49",
X"E13D",
X"D48B",
X"D96D",
X"D314",
X"D48B",
X"D314",
X"DA67",
X"D314",
X"CF2C",
X"D9EA",
X"DAE4",
X"D67F",
X"D48B",
X"DCD8",
X"DB61",
X"D6FC",
X"D96D",
X"E0C0",
X"D8F0",
X"D8F0",
X"D9EA",
X"D96D",
X"DE4F",
X"E043",
X"EE6C",
X"DF49",
X"EFE3",
X"F4C5",
X"F92A",
X"07D0",
X"FF83",
X"0BB8",
X"128E",
X"1405",
X"1B58",
X"2599",
X"1B58",
X"2710",
X"2616",
X"2FDA",
X"2E63",
X"2422",
X"278D",
X"2981",
X"3151",
X"203A",
X"2904",
X"2887",
X"203A",
X"2328",
X"203A",
X"29FE",
X"222E",
X"2D69",
X"29FE",
X"2710",
X"2710",
X"2B75",
X"2E63",
X"2710",
X"21B1",
X"1C52",
X"20B7",
X"1F40",
X"2616",
X"19E1",
X"15F9",
X"0FA0",
X"1405",
X"08CA",
X"08CA",
X"04E2",
X"F7B3",
X"F34E",
X"E61F",
X"EB01",
X"E237",
X"DBDE",
X"DCD8",
X"DA67",
X"D391",
X"DAE4",
X"E043",
X"D7F6",
X"DC5B",
X"E13D",
X"D6FC",
X"EDEF",
X"E42B",
X"E813",
X"EA07",
X"F2D1",
X"FE89",
X"F830",
X"05DC",
X"F9A7",
X"0753",
X"0ABE",
X"084D",
X"1388",
X"036B",
X"0D2F",
X"0ABE",
X"0C35",
X"0CB2",
X"0FA0",
X"101D",
X"128E",
X"0659",
X"FD12",
X"F8AD",
X"ECF5",
X"F15A",
X"DBDE",
X"E237",
X"DE4F",
X"DF49",
X"DF49",
X"D21A",
X"DE4F",
X"D6FC",
X"E890",
X"D508",
X"E0C0",
X"D873",
X"DE4F",
X"E98A",
X"DECC",
X"F15A",
X"E5A2",
X"F7B3",
X"F060",
X"007D",
X"F34E",
X"FD8F",
X"0BB8",
X"0177",
X"0659",
X"0271",
X"0177",
X"F63C",
X"FD12",
X"F5BF",
X"FF06",
X"FF83",
X"02EE",
X"109A",
X"07D0",
X"1405",
X"1CCF",
X"1FBD",
X"1E46",
X"21B1",
X"2CEC",
X"2328",
X"251C",
X"2D69",
X"21B1",
X"20B7",
X"2A7B",
X"278D",
X"1B58",
X"130B",
X"2616",
X"1BD5",
X"1EC3",
X"2E63",
X"2887",
X"1CCF",
X"2A7B",
X"1EC3",
X"1770",
X"1BD5",
X"1FBD",
X"16F3",
X"109A",
X"2599",
X"280A",
X"19E1",
X"2AF8",
X"2134",
X"1DC9",
X"2616",
X"1F40",
X"29FE",
X"14FF",
X"186A",
X"203A",
X"1BD5",
X"21B1",
X"22AB",
X"1FBD",
X"1482",
X"084D",
X"FD8F",
X"F9A7",
X"F92A",
X"F254",
X"F9A7",
X"F63C",
X"EB01",
X"F6B9",
X"EF66",
X"F254",
X"F1D7",
X"F2D1",
X"F15A",
X"FD8F",
X"F7B3",
X"04E2",
X"0000",
X"084D",
X"0947",
X"0947",
X"1ADB",
X"01F4",
X"16F3",
X"157C",
X"1E46",
X"1A5E",
X"22AB",
X"19E1",
X"1388",
X"203A",
X"1388",
X"109A",
X"1194",
X"0F23",
X"0C35",
X"0947",
X"0A41",
X"00FA",
X"F9A7",
X"F8AD",
X"F92A",
X"EA07",
X"FD12",
X"EF66",
X"F254",
X"F6B9",
X"EF66",
X"F7B3",
X"EBFB",
X"F254",
X"F92A",
X"EF66",
X"F2D1",
X"F0DD",
X"EFE3",
X"EC78",
X"EB01",
X"EC78",
X"EBFB",
X"E525",
X"DBDE",
X"E1BA",
X"DECC",
X"DA67",
X"D508",
X"DF49",
X"D9EA",
X"D602",
X"E0C0",
X"D9EA",
X"E331",
X"E0C0",
X"E3AE",
X"E90D",
X"E1BA",
X"E90D",
X"F15A",
X"EE6C",
X"E61F",
X"F15A",
X"EE6C",
X"ECF5",
X"ECF5",
X"F15A",
X"EB01",
X"F254",
X"E813",
X"EB01",
X"E525",
X"E69C",
X"E5A2",
X"E5A2",
X"E796",
X"DCD8",
X"E2B4",
X"E331",
X"DA67",
X"DFC6",
X"DECC",
X"CFA9",
X"E237",
X"DCD8",
X"D602",
X"DF49",
X"D508",
X"E331",
X"DB61",
X"DFC6",
X"E42B",
X"E043",
X"DC5B",
X"F0DD",
X"E796",
X"DDD2",
X"F6B9",
X"F1D7",
X"EE6C",
X"FD12",
X"F63C",
X"F830",
X"0753",
X"F8AD",
X"03E8",
X"05DC",
X"F9A7",
X"07D0",
X"FAA1",
X"0753",
X"09C4",
X"0753",
X"0F23",
X"09C4",
X"1194",
X"1964",
X"157C",
X"186A",
X"1194",
X"130B",
X"1388",
X"0FA0",
X"02EE",
X"FD12",
X"F92A",
X"EBFB",
X"E796",
X"E69C",
X"F2D1",
X"F8AD",
X"05DC",
X"02EE",
X"0659",
X"F542",
X"0000",
X"FB9B",
X"F830",
X"FD8F",
X"F63C",
X"F7B3",
X"FC18",
X"FB9B",
X"F8AD",
X"05DC",
X"00FA",
X"F7B3",
X"0000",
X"036B",
X"FE0C",
X"FF06",
X"0000",
X"09C4",
X"15F9",
X"1117",
X"130B",
X"14FF",
X"09C4",
X"007D",
X"03E8",
X"EBFB",
X"EF66",
X"F3CB",
X"F448",
X"FB1E",
X"09C4",
X"0177",
X"07D0",
X"0F23",
X"0465",
X"055F",
X"1194",
X"1211",
X"0465",
X"1388",
X"222E",
X"1CCF",
X"2BF2",
X"2FDA",
X"2616",
X"3057",
X"2E63",
X"1A5E",
X"1ADB",
X"1388",
X"15F9",
X"17ED",
X"186A",
X"17ED",
X"21B1",
X"2422",
X"2904",
X"2CEC",
X"2CEC",
X"2AF8",
X"249F",
X"29FE",
X"2710",
X"2BF2",
X"23A5",
X"249F",
X"1FBD",
X"22AB",
X"249F",
X"2DE6",
X"2C6F",
X"2AF8",
X"2BF2",
X"2904",
X"21B1",
X"1DC9",
X"22AB",
X"21B1",
X"20B7",
X"1F40",
X"1ADB",
X"1BD5",
X"1482",
X"1211",
X"14FF",
X"0B3B",
X"0F23",
X"101D",
X"02EE",
X"0271",
X"00FA",
X"FC18",
X"FC18",
X"F3CB",
X"F060",
X"F254",
X"F736",
X"E890",
X"F5BF",
X"E890",
X"EA07",
X"E98A",
X"D873",
X"D602",
X"D0A3",
X"DC5B",
X"D602",
X"D7F6",
X"EB01",
X"DF49",
X"E043",
X"DAE4",
X"DECC",
X"CDB5",
X"CE32",
X"D40E",
X"CEAF",
X"D6FC",
X"D779",
X"D19D",
X"D297",
X"DD55",
X"DC5B",
X"D508",
X"D40E",
X"DC5B",
X"D120",
X"DC5B",
X"D48B",
X"DA67",
X"D8F0",
X"DBDE",
X"E796",
X"E331",
X"DFC6",
X"E2B4",
X"DD55",
X"E5A2",
X"E61F",
X"F060",
X"ECF5",
X"EF66",
X"FB1E",
X"F254",
X"F9A7",
X"F254",
X"00FA",
X"F448",
X"0271",
X"FF06",
X"F830",
X"F9A7",
X"F9A7",
X"F736",
X"F542",
X"F448",
X"ED72",
X"F0DD",
X"F254",
X"EF66",
X"F1D7",
X"F15A",
X"F15A",
X"F9A7",
X"F92A",
X"F9A7",
X"F830",
X"0753",
X"FC95",
X"FB9B",
X"0271",
X"F92A",
X"02EE",
X"F9A7",
X"1117",
X"FA24",
X"0753",
X"FB1E",
X"01F4",
X"0177",
X"01F4",
X"08CA",
X"06D6",
X"0F23",
X"0ABE",
X"1F40",
X"1ADB",
X"130B",
X"222E",
X"18E7",
X"19E1",
X"084D",
X"14FF",
X"186A",
X"0F23",
X"128E",
X"0B3B",
X"0E29",
X"FAA1",
X"F9A7",
X"FD12",
X"F6B9",
X"F2D1",
X"F060",
X"02EE",
X"FC95",
X"0ABE",
X"0CB2",
X"0CB2",
X"0D2F",
X"0ABE",
X"09C4",
X"00FA",
X"0ABE",
X"0EA6",
X"055F",
X"14FF",
X"186A",
X"2887",
X"29FE",
X"22AB",
X"31CE",
X"3345",
X"2DE6",
X"2E63",
X"2E63",
X"2904",
X"186A",
X"130B",
X"2887",
X"0E29",
X"1A5E",
X"1CCF",
X"1C52",
X"22AB",
X"21B1",
X"21B1",
X"2328",
X"2B75",
X"2693",
X"2981",
X"2D69",
X"1EC3",
X"2422",
X"249F",
X"2887",
X"2E63",
X"2328",
X"20B7",
X"203A",
X"15F9",
X"1B58",
X"186A",
X"1B58",
X"1482",
X"1EC3",
X"2328",
X"17ED",
X"1DC9",
X"21B1",
X"15F9",
X"1CCF",
X"2599",
X"1B58",
X"2134",
X"2328",
X"2693",
X"1FBD",
X"1A5E",
X"1F40",
X"0CB2",
X"1388",
X"09C4",
X"FC18",
X"0177",
X"FD8F",
X"F448",
X"EBFB",
X"EBFB",
X"E4A8",
X"EEE9",
X"E237",
X"DC5B",
X"D602",
X"DF49",
X"D779",
X"DB61",
X"DE4F",
X"E237",
X"D7F6",
X"CD38",
X"D7F6",
X"D391",
X"D391",
X"DAE4",
X"D8F0",
X"F1D7",
X"DD55",
X"E719",
X"EDEF",
X"DFC6",
X"DE4F",
X"DAE4",
X"D602",
X"DC5B",
X"D873",
X"DFC6",
X"DCD8",
X"DD55",
X"DCD8",
X"D873",
X"DC5B",
X"D297",
X"DB61",
X"D585",
X"CEAF",
X"D602",
X"CC3E",
X"DAE4",
X"D7F6",
X"DB61",
X"DE4F",
X"E13D",
X"E1BA",
X"F0DD",
X"0177",
X"FE89",
X"F9A7",
X"036B",
X"0DAC",
X"FF06",
X"0177",
X"FF83",
X"0659",
X"F830",
X"F542",
X"EEE9",
X"F0DD",
X"F448",
X"EA84",
X"EE6C",
X"E043",
X"E0C0",
X"D6FC",
X"D585",
X"D026",
X"D873",
X"D602",
X"DAE4",
X"DE4F",
X"D96D",
X"DECC",
X"E4A8",
X"E69C",
X"E42B",
X"F060",
X"F6B9",
X"ED72",
X"FA24",
X"F9A7",
X"055F",
X"08CA",
X"0BB8",
X"0EA6",
X"0FA0",
X"186A",
X"1482",
X"17ED",
X"1211",
X"1CCF",
X"186A",
X"186A",
X"17ED",
X"1ADB",
X"1B58",
X"1BD5",
X"101D",
X"109A",
X"1B58",
X"1964",
X"2134",
X"1EC3",
X"1FBD",
X"2134",
X"1B58",
X"1ADB",
X"1ADB",
X"1CCF",
X"1A5E",
X"1964",
X"186A",
X"1676",
X"1770",
X"1211",
X"1194",
X"0E29",
X"084D",
X"00FA",
X"02EE",
X"0A41",
X"01F4",
X"01F4",
X"0ABE",
X"14FF",
X"17ED",
X"1770",
X"1676",
X"1482",
X"18E7",
X"1A5E",
X"1B58",
X"222E",
X"251C",
X"222E",
X"23A5",
X"2599",
X"2F5D",
X"2D69",
X"2A7B",
X"2A7B",
X"2616",
X"2C6F",
X"2422",
X"2134",
X"2599",
X"1F40",
X"1FBD",
X"1FBD",
X"186A",
X"0CB2",
X"0DAC",
X"1211",
X"0465",
X"0BB8",
X"128E",
X"09C4",
X"0B3B",
X"0DAC",
X"0A41",
X"0EA6",
X"036B",
X"FD12",
X"F7B3",
X"EFE3",
X"EB01",
X"EC78",
X"E1BA",
X"F5BF",
X"EFE3",
X"F060",
X"FA24",
X"007D",
X"0271",
X"F9A7",
X"FE0C",
X"0271",
X"F8AD",
X"01F4",
X"FE0C",
X"F92A",
X"0A41",
X"FB9B",
X"FB9B",
X"F8AD",
X"FE89",
X"FC18",
X"F9A7",
X"FB9B",
X"FAA1",
X"EA84",
X"EA07",
X"E796",
X"E525",
X"ED72",
X"E525",
X"D96D",
X"E719",
X"DC5B",
X"DECC",
X"D873",
X"DB61",
X"DF49",
X"DA67",
X"DA67",
X"D120",
X"E3AE",
X"CF2C",
X"DA67",
X"D7F6",
X"D9EA",
X"DD55",
X"D585",
X"DDD2",
X"E237",
X"ECF5",
X"E5A2",
X"DECC",
X"EC78",
X"EE6C",
X"EEE9",
X"F254",
X"F830",
X"F2D1",
X"F2D1",
X"FA24",
X"F3CB",
X"00FA",
X"0465",
X"F34E",
X"F448",
X"F448",
X"F542",
X"F5BF",
X"EC78",
X"F3CB",
X"E90D",
X"F542",
X"E90D",
X"F4C5",
X"F92A",
X"F542",
X"F1D7",
X"F254",
X"EF66",
X"F4C5",
X"01F4",
X"F1D7",
X"0000",
X"F830",
X"F7B3",
X"F3CB",
X"F6B9",
X"0947",
X"055F",
X"02EE",
X"0177",
X"FAA1",
X"FD12",
X"F63C",
X"F8AD",
X"F830",
X"FE89",
X"0271",
X"FD8F",
X"055F",
X"0BB8",
X"1211",
X"15F9",
X"1D4C",
X"251C",
X"1E46",
X"203A",
X"251C",
X"2616",
X"1FBD",
X"1CCF",
X"19E1",
X"0D2F",
X"1117",
X"0CB2",
X"07D0",
X"0659",
X"FF06",
X"FF06",
X"0177",
X"F92A",
X"FB1E",
X"F63C",
X"F9A7",
X"F6B9",
X"F92A",
X"F63C",
X"F736",
X"FC18",
X"F8AD",
X"F3CB",
X"F9A7",
X"FA24",
X"F448",
X"007D",
X"FC18",
X"F4C5",
X"FB9B",
X"FE0C",
X"F6B9",
X"FE89",
X"F830",
X"FB9B",
X"F1D7",
X"F542",
X"FA24",
X"0465",
X"084D",
X"FE0C",
X"06D6",
X"055F",
X"FB9B",
X"03E8",
X"0C35",
X"04E2",
X"0A41",
X"04E2",
X"0ABE",
X"18E7",
X"1211",
X"186A",
X"203A",
X"1BD5",
X"1C52",
X"1CCF",
X"1EC3",
X"1C52",
X"2599",
X"1CCF",
X"1CCF",
X"22AB",
X"1DC9",
X"278D",
X"2134",
X"22AB",
X"2B75",
X"2904",
X"2AF8",
X"2422",
X"2904",
X"2AF8",
X"29FE",
X"280A",
X"2328",
X"2A7B",
X"2599",
X"2710",
X"1EC3",
X"1770",
X"1F40",
X"1C52",
X"1FBD",
X"1DC9",
X"17ED",
X"1A5E",
X"17ED",
X"1388",
X"1117",
X"0DAC",
X"0ABE",
X"FD12",
X"FF83",
X"F830",
X"02EE",
X"FE0C",
X"06D6",
X"0271",
X"FF06",
X"0177",
X"FF06",
X"0753",
X"05DC",
X"FD8F",
X"0271",
X"0271",
X"FAA1",
X"FD8F",
X"FE89",
X"0271",
X"FC18",
X"F8AD",
X"0753",
X"03E8",
X"F736",
X"0465",
X"0000",
X"FC18",
X"F542",
X"FE89",
X"FE89",
X"F736",
X"F8AD",
X"F448",
X"F448",
X"E890",
X"ED72",
X"E813",
X"DC5B",
X"D96D",
X"DDD2",
X"DCD8",
X"D779",
X"D779",
X"D779",
X"D779",
X"D19D",
X"D7F6",
X"D40E",
X"DBDE",
X"D96D",
X"DC5B",
X"DECC",
X"E043",
X"E0C0",
X"EA07",
X"EB7E",
X"E719",
X"ED72",
X"F060",
X"F5BF",
X"ECF5",
X"EA84",
X"F060",
X"F15A",
X"F4C5",
X"F2D1",
X"FB1E",
X"FE0C",
X"FC18",
X"03E8",
X"04E2",
X"FE89",
X"036B",
X"055F",
X"0177",
X"03E8",
X"FC18",
X"F736",
X"FA24",
X"F8AD",
X"F6B9",
X"FB1E",
X"F34E",
X"FAA1",
X"F830",
X"F6B9",
X"F9A7",
X"F34E",
X"F8AD",
X"FAA1",
X"FD8F",
X"F92A",
X"FAA1",
X"F830",
X"F8AD",
X"F9A7",
X"F63C",
X"F8AD",
X"F4C5",
X"F4C5",
X"F542",
X"F060",
X"F15A",
X"F1D7",
X"F1D7",
X"F0DD",
X"EF66",
X"F15A",
X"E525",
X"E61F",
X"E69C",
X"E98A",
X"E525",
X"DC5B",
X"E69C",
X"E813",
X"EDEF",
X"F254",
X"F1D7",
X"F4C5",
X"F736",
X"FAA1",
X"FF83",
X"007D",
X"0947",
X"0A41",
X"0E29",
X"128E",
X"15F9",
X"1770",
X"16F3",
X"186A",
X"1D4C",
X"1BD5",
X"1D4C",
X"2422",
X"2422",
X"278D",
X"23A5",
X"2D69",
X"280A",
X"278D",
X"2422",
X"23A5",
X"249F",
X"2981",
X"2599",
X"2710",
X"2616",
X"1CCF",
X"1ADB",
X"1C52",
X"1FBD",
X"1194",
X"1676",
X"0F23",
X"0E29",
X"1117",
X"0947",
X"0ABE",
X"04E2",
X"FF83",
X"FD8F",
X"F9A7",
X"F2D1",
X"F254",
X"ED72",
X"E237",
X"E0C0",
X"E1BA",
X"DD55",
X"D8F0",
X"DECC",
X"D8F0",
X"D873",
X"D779",
X"D7F6",
X"D873",
X"D6FC",
X"E1BA",
X"E1BA",
X"E42B",
X"E237",
X"EE6C",
X"F15A",
X"F448",
X"F63C",
X"F542",
X"FC95",
X"FAA1",
X"0465",
X"FE89",
X"055F",
X"0465",
X"F63C",
X"FAA1",
X"0000",
X"FF83",
X"06D6",
X"0000",
X"036B",
X"0753",
X"FF83",
X"0B3B",
X"FF06",
X"FF06",
X"08CA",
X"0659",
X"08CA",
X"00FA",
X"0659",
X"007D",
X"02EE",
X"0465",
X"F9A7",
X"FD12",
X"F736",
X"F830",
X"F448",
X"FAA1",
X"F92A",
X"FF06",
X"FE89",
X"04E2",
X"0ABE",
X"02EE",
X"0D2F",
X"0C35",
X"0753",
X"07D0",
X"0CB2",
X"0947",
X"09C4",
X"0BB8",
X"109A",
X"0D2F",
X"0A41",
X"0ABE",
X"0CB2",
X"084D",
X"05DC",
X"03E8",
X"04E2",
X"0465",
X"FD12",
X"0271",
X"FE89",
X"FAA1",
X"F92A",
X"F830",
X"F8AD",
X"F060",
X"F6B9",
X"F736",
X"EB01",
X"ECF5",
X"E61F",
X"E331",
X"E42B",
X"DE4F",
X"D9EA",
X"E2B4",
X"DD55",
X"DFC6",
X"E237",
X"E043",
X"D8F0",
X"E0C0",
X"E331",
X"DB61",
X"E90D",
X"DF49",
X"E69C",
X"E42B",
X"E237",
X"EDEF",
X"E890",
X"EEE9",
X"F448",
X"FC95",
X"FD12",
X"F7B3",
X"00FA",
X"03E8",
X"0753",
X"0947",
X"08CA",
X"0E29",
X"0EA6",
X"0DAC",
X"0CB2",
X"0E29",
X"0C35",
X"0EA6",
X"0C35",
X"0B3B",
X"0ABE",
X"1117",
X"0C35",
X"1676",
X"0659",
X"08CA",
X"1770",
X"0F23",
X"1E46",
X"20B7",
X"1FBD",
X"1676",
X"17ED",
X"1A5E",
X"1405",
X"186A",
X"1482",
X"1A5E",
X"203A",
X"15F9",
X"1F40",
X"1E46",
X"2134",
X"2710",
X"21B1",
X"1CCF",
X"21B1",
X"1C52",
X"2887",
X"1CCF",
X"16F3",
X"1DC9",
X"18E7",
X"222E",
X"1C52",
X"1A5E",
X"16F3",
X"14FF",
X"1770",
X"1388",
X"17ED",
X"1B58",
X"1C52",
X"2328",
X"251C",
X"2887",
X"23A5",
X"2328",
X"222E",
X"2134",
X"2599",
X"1B58",
X"2693",
X"1EC3",
X"249F",
X"2134",
X"222E",
X"2599",
X"23A5",
X"278D",
X"203A",
X"2693",
X"22AB",
X"203A",
X"1C52",
X"1ADB",
X"1770",
X"17ED",
X"109A",
X"16F3",
X"1C52",
X"128E",
X"186A",
X"1194",
X"1211",
X"1482",
X"0C35",
X"0D2F",
X"0C35",
X"0465",
X"0C35",
X"FF06",
X"02EE",
X"07D0",
X"03E8",
X"0659",
X"06D6",
X"03E8",
X"04E2",
X"0ABE",
X"101D",
X"0CB2",
X"0F23",
X"130B",
X"0B3B",
X"0F23",
X"1482",
X"130B",
X"084D",
X"130B",
X"1194",
X"19E1",
X"1211",
X"101D",
X"0F23",
X"03E8",
X"07D0",
X"FC95",
X"FF06",
X"F34E",
X"F92A",
X"F254",
X"E796",
X"E69C",
X"DCD8",
X"DBDE",
X"D602",
X"D6FC",
X"D7F6",
X"DA67",
X"D67F",
X"D8F0",
X"D873",
X"D48B",
X"D9EA",
X"CDB5",
X"CE32",
X"D19D",
X"CD38",
X"D21A",
X"C950",
X"CE32",
X"D48B",
X"CF2C",
X"D026",
X"CF2C",
X"CDB5",
X"C950",
X"CE32",
X"D120",
X"CD38",
X"CB44",
X"CDB5",
X"D0A3",
X"CD38",
X"CD38",
X"CBC1",
X"D0A3",
X"CCBB",
X"CD38",
X"CDB5",
X"C8D3",
X"CEAF",
X"C9CD",
X"D120",
X"D120",
X"D508",
X"D120",
X"D40E",
X"D67F",
X"D508",
X"D602",
X"D602",
X"D602",
X"D873",
X"D585",
X"D96D",
X"DBDE",
X"DA67",
X"DCD8",
X"DDD2",
X"DF49",
X"D7F6",
X"DCD8",
X"DAE4",
X"DE4F",
X"E525",
X"D9EA",
X"E796",
X"E90D",
X"EB7E",
X"F15A",
X"EA84",
X"F4C5",
X"F448",
X"F4C5",
X"FB1E",
X"FD8F",
X"FF83",
X"FD8F",
X"0465",
X"0B3B",
X"0753",
X"09C4",
X"0C35",
X"0A41",
X"1117",
X"109A",
X"15F9",
X"1676",
X"157C",
X"2328",
X"1E46",
X"1EC3",
X"2134",
X"2328",
X"2904",
X"23A5",
X"21B1",
X"30D4",
X"251C",
X"3057",
X"3057",
X"2BF2",
X"2BF2",
X"2E63",
X"33C2",
X"2D69",
X"32C8",
X"31CE",
X"2887",
X"2FDA",
X"34BC",
X"2693",
X"34BC",
X"2BF2",
X"2B75",
X"3151",
X"2FDA",
X"35B6",
X"2FDA",
X"2CEC",
X"324B",
X"2BF2",
X"2FDA",
X"2BF2",
X"2E63",
X"2FDA",
X"2693",
X"32C8",
X"2887",
X"29FE",
X"280A",
X"2904",
X"23A5",
X"280A",
X"2599",
X"20B7",
X"2422",
X"20B7",
X"2BF2",
X"23A5",
X"1DC9",
X"2981",
X"22AB",
X"1BD5",
X"29FE",
X"1F40",
X"1FBD",
X"2599",
X"23A5",
X"2616",
X"249F",
X"2BF2",
X"2710",
X"23A5",
X"2693",
X"249F",
X"23A5",
X"2134",
X"2599",
X"1E46",
X"1E46",
X"1FBD",
X"1A5E",
X"19E1",
X"1ADB",
X"109A",
X"0EA6",
X"0271",
X"FC18",
X"F92A",
X"F92A",
X"F15A",
X"F448",
X"FB1E",
X"F6B9",
X"F5BF",
X"FC95",
X"FC18",
X"F736",
X"EE6C",
X"F15A",
X"EB7E",
X"E796",
X"EC78",
X"E3AE",
X"DD55",
X"DECC",
X"E0C0",
X"D6FC",
X"DB61",
X"D19D",
X"D120",
X"D297",
X"CBC1",
X"D026",
X"D120",
X"CDB5",
X"C9CD",
X"D026",
X"CFA9",
X"C5E5",
X"C662",
X"C374",
X"CDB5",
X"CA4A",
X"CDB5",
X"C9CD",
X"D0A3",
X"D873",
X"D21A",
X"D40E",
X"D48B",
X"D7F6",
X"D21A",
X"D779",
X"D297",
X"D026",
X"CD38",
X"CE32",
X"D48B",
X"D026",
X"D026",
X"D67F",
X"D9EA",
X"D6FC",
X"D779",
X"DBDE",
X"DC5B",
X"DD55",
X"DE4F",
X"E0C0",
X"E525",
X"E13D",
X"E796",
X"EDEF",
X"F448",
X"EEE9",
X"F5BF",
X"FF83",
X"FAA1",
X"01F4",
X"02EE",
X"FD12",
X"0A41",
X"03E8",
X"036B",
X"0B3B",
X"0753",
X"055F",
X"0C35",
X"0CB2",
X"FF06",
X"00FA",
X"0E29",
X"0271",
X"036B",
X"0B3B",
X"FE89",
X"0659",
X"07D0",
X"0465",
X"02EE",
X"0659",
X"02EE",
X"03E8",
X"0271",
X"05DC",
X"0F23",
X"0C35",
X"0A41",
X"08CA",
X"0A41",
X"01F4",
X"0BB8",
X"0000",
X"07D0",
X"036B",
X"0177",
X"0EA6",
X"0BB8",
X"055F",
X"1482",
X"0D2F",
X"0E29",
X"157C",
X"1770",
X"0EA6",
X"0FA0",
X"1117",
X"101D",
X"08CA",
X"06D6",
X"0B3B",
X"08CA",
X"084D",
X"06D6",
X"0ABE",
X"0C35",
X"0271",
X"09C4",
X"0659",
X"0ABE",
X"08CA",
X"0947",
X"08CA",
X"0465",
X"0DAC",
X"0BB8",
X"0A41",
X"0CB2",
X"0947",
X"0EA6",
X"157C",
X"1EC3",
X"2422",
X"1DC9",
X"1D4C",
X"2AF8",
X"2710",
X"2B75",
X"249F",
X"2693",
X"280A",
X"1FBD",
X"1F40",
X"1B58",
X"18E7",
X"186A",
X"1DC9",
X"2134",
X"1BD5",
X"1B58",
X"22AB",
X"1C52",
X"1676",
X"1482",
X"16F3",
X"130B",
X"0ABE",
X"1482",
X"0FA0",
X"0FA0",
X"101D",
X"128E",
X"14FF",
X"1405",
X"1405",
X"1194",
X"1676",
X"1405",
X"15F9",
X"19E1",
X"1676",
X"1964",
X"249F",
X"2616",
X"2616",
X"21B1",
X"2328",
X"2693",
X"1DC9",
X"1FBD",
X"2328",
X"1EC3",
X"1F40",
X"222E",
X"1ADB",
X"1C52",
X"1A5E",
X"1770",
X"17ED",
X"157C",
X"1194",
X"0F23",
X"0EA6",
X"0A41",
X"05DC",
X"0C35",
X"07D0",
X"0BB8",
X"04E2",
X"0DAC",
X"0465",
X"0753",
X"0A41",
X"0271",
X"09C4",
X"F9A7",
X"FAA1",
X"036B",
X"F8AD",
X"01F4",
X"F6B9",
X"F6B9",
X"F34E",
X"ECF5",
X"EEE9",
X"E61F",
X"E5A2",
X"DE4F",
X"E61F",
X"E2B4",
X"E1BA",
X"E813",
X"E69C",
X"E719",
X"DCD8",
X"E5A2",
X"E1BA",
X"E796",
X"E13D",
X"E69C",
X"E796",
X"E2B4",
X"E525",
X"E3AE",
X"D9EA",
X"DD55",
X"D6FC",
X"D19D",
X"CEAF",
X"D21A",
X"CCBB",
X"CCBB",
X"D026",
X"CAC7",
X"D297",
X"CB44",
X"D19D",
X"CC3E",
X"D026",
X"CC3E",
X"D120",
X"D0A3",
X"CB44",
X"CD38",
X"D21A",
X"D19D",
X"CCBB",
X"D21A",
X"D0A3",
X"CAC7",
X"CDB5",
X"CE32",
X"CEAF",
X"CFA9",
X"D026",
X"D297",
X"CE32",
X"D48B",
X"D314",
X"DA67",
X"D21A",
X"D9EA",
X"D9EA",
X"D391",
X"DECC",
X"D8F0",
X"DECC",
X"E0C0",
X"E331",
X"DB61",
X"DFC6",
X"DC5B",
X"E043",
X"E42B",
X"DAE4",
X"E237",
X"E525",
X"E61F",
X"DD55",
X"E42B",
X"E61F",
X"EB7E",
X"E61F",
X"EA84",
X"E813",
X"F63C",
X"ED72",
X"F448",
X"F736",
X"F254",
X"F7B3",
X"F7B3",
X"FD12",
X"FA24",
X"FAA1",
X"FB9B",
X"FB1E",
X"FC18",
X"FAA1",
X"FE89",
X"007D",
X"04E2",
X"05DC",
X"07D0",
X"1117",
X"1211",
X"14FF",
X"1388",
X"157C",
X"1B58",
X"1964",
X"1CCF",
X"2134",
X"20B7",
X"280A",
X"280A",
X"2AF8",
X"2AF8",
X"2904",
X"2422",
X"2904",
X"2328",
X"2693",
X"222E",
X"2A7B",
X"2A7B",
X"2D69",
X"2D69",
X"2CEC",
X"31CE",
X"3345",
X"34BC",
X"2F5D",
X"36B0",
X"33C2",
X"324B",
X"3539",
X"3539",
X"343F",
X"343F",
X"35B6",
X"34BC",
X"3633",
X"3539",
X"34BC",
X"3151",
X"2FDA",
X"2EE0",
X"2DE6",
X"2E63",
X"30D4",
X"2BF2",
X"2AF8",
X"2D69",
X"2CEC",
X"2F5D",
X"2981",
X"2EE0",
X"2AF8",
X"2C6F",
X"2887",
X"2AF8",
X"278D",
X"2693",
X"280A",
X"2422",
X"249F",
X"2328",
X"22AB",
X"1EC3",
X"21B1",
X"1A5E",
X"18E7",
X"186A",
X"1388",
X"14FF",
X"0D2F",
X"0BB8",
X"0A41",
X"02EE",
X"00FA",
X"06D6",
X"03E8",
X"00FA",
X"00FA",
X"007D",
X"FE0C",
X"FB1E",
X"F448",
X"F0DD",
X"ED72",
X"E90D",
X"EA07",
X"E69C",
X"EA84",
X"E890",
X"E90D",
X"E525",
X"E3AE",
X"DBDE",
X"DB61",
X"D297",
X"D6FC",
X"D314",
X"CF2C",
X"D314",
X"C662",
X"C5E5",
X"C662",
X"C4EB",
X"C856",
X"C3F1",
X"C9CD",
X"C6DF",
X"C8D3",
X"CB44",
X"CF2C",
X"D120",
X"D0A3",
X"D508",
X"D21A",
X"D67F",
X"CFA9",
X"D67F",
X"DA67",
X"D67F",
X"D585",
X"D7F6",
X"DF49",
X"E4A8",
X"E0C0",
X"DF49",
X"F060",
X"E813",
X"E61F",
X"ED72",
X"ED72",
X"EF66",
X"F15A",
X"F6B9",
X"F8AD",
X"FA24",
X"F6B9",
X"F2D1",
X"EF66",
X"E5A2",
X"EA84",
X"EEE9",
X"E331",
X"E13D",
X"ECF5",
X"EA07",
X"E69C",
X"EEE9",
X"E719",
X"E98A",
X"F3CB",
X"E890",
X"EEE9",
X"EF66",
X"E61F",
X"EE6C",
X"F542",
X"EF66",
X"F448",
X"F254",
X"F34E",
X"F4C5",
X"F830",
X"F34E",
X"EFE3",
X"FAA1",
X"F15A",
X"F7B3",
X"F830",
X"F3CB",
X"F8AD",
X"FD8F",
X"FAA1",
X"00FA",
X"F830",
X"FC95",
X"02EE",
X"F542",
X"036B",
X"FE89",
X"0000",
X"0753",
X"FF06",
X"05DC",
X"05DC",
X"FC95",
X"0BB8",
X"FD12",
X"04E2",
X"0271",
X"0659",
X"02EE",
X"06D6",
X"0ABE",
X"0465",
X"130B",
X"0C35",
X"05DC",
X"157C",
X"1194",
X"1BD5",
X"1482",
X"17ED",
X"1CCF",
X"1B58",
X"1770",
X"14FF",
X"1CCF",
X"0CB2",
X"1BD5",
X"15F9",
X"2134",
X"19E1",
X"2422",
X"249F",
X"1FBD",
X"22AB",
X"2C6F",
X"2616",
X"2599",
X"32C8",
X"22AB",
X"2EE0",
X"3057",
X"2AF8",
X"38A4",
X"324B",
X"2B75",
X"3539",
X"2B75",
X"2904",
X"2328",
X"22AB",
X"2887",
X"278D",
X"2887",
X"2904",
X"278D",
X"1DC9",
X"249F",
X"1B58",
X"157C",
X"1117",
X"1405",
X"1ADB",
X"1EC3",
X"2616",
X"2710",
X"2710",
X"23A5",
X"2134",
X"222E",
X"0D2F",
X"1676",
X"1F40",
X"0EA6",
X"084D",
X"1117",
X"084D",
X"02EE",
X"1405",
X"0D2F",
X"055F",
X"0271",
X"FD12",
X"FD12",
X"F542",
X"EBFB",
X"EF66",
X"EE6C",
X"F060",
X"EDEF",
X"EA07",
X"E813",
X"EB01",
X"E42B",
X"E043",
X"E13D",
X"DC5B",
X"D96D",
X"DD55",
X"D0A3",
X"D314",
X"D21A",
X"D21A",
X"D0A3",
X"C950",
X"CA4A",
X"CB44",
X"CE32",
X"CA4A",
X"CC3E",
X"C856",
X"C950",
X"C8D3",
X"C8D3",
X"C950",
X"C950",
X"C9CD",
X"D19D",
X"D40E",
X"D6FC",
X"D8F0",
X"D7F6",
X"D8F0",
X"DBDE",
X"D297",
X"D0A3",
X"D391",
X"CE32",
X"D67F",
X"D585",
X"D508",
X"D8F0",
X"DDD2",
X"D8F0",
X"D6FC",
X"D19D",
X"D602",
X"D779",
X"D67F",
X"D6FC",
X"D96D",
X"D96D",
X"E61F",
X"DFC6",
X"E0C0",
X"E98A",
X"E3AE",
X"E61F",
X"F3CB",
X"F542",
X"F1D7",
X"FC18",
X"01F4",
X"01F4",
X"0177",
X"03E8",
X"0C35",
X"1482",
X"157C",
X"1405",
X"1770",
X"1117",
X"101D",
X"1DC9",
X"1D4C",
X"1F40",
X"1DC9",
X"1F40",
X"249F",
X"2887",
X"2710",
X"2134",
X"2134",
X"15F9",
X"18E7",
X"1ADB",
X"1DC9",
X"1FBD",
X"2134",
X"1FBD",
X"20B7",
X"2599",
X"2599",
X"2BF2",
X"2887",
X"3151",
X"2A7B",
X"2A7B",
X"3539",
X"2904",
X"34BC",
X"343F",
X"2D69",
X"3539",
X"2FDA",
X"2EE0",
X"31CE",
X"31CE",
X"2E63",
X"2B75",
X"280A",
X"249F",
X"2328",
X"222E",
X"1DC9",
X"1C52",
X"1DC9",
X"1A5E",
X"1964",
X"1A5E",
X"157C",
X"1964",
X"1405",
X"0C35",
X"05DC",
X"08CA",
X"0B3B",
X"0271",
X"0177",
X"09C4",
X"0000",
X"05DC",
X"FF06",
X"F830",
X"036B",
X"F9A7",
X"F5BF",
X"F254",
X"ED72",
X"EE6C",
X"E69C",
X"E796",
X"E3AE",
X"E69C",
X"E90D",
X"E813",
X"E890",
X"E525",
X"E5A2",
X"EA07",
X"E043",
X"E4A8",
X"E90D",
X"E043",
X"E3AE",
X"E5A2",
X"E890",
X"E42B",
X"E237",
X"E1BA",
X"E42B",
X"E61F",
X"E5A2",
X"EC78",
X"E796",
X"E890",
X"ECF5",
X"EDEF",
X"EA07",
X"EBFB",
X"EE6C",
X"EBFB",
X"ECF5",
X"F15A",
X"F060",
X"EA84",
X"EA84",
X"EB7E",
X"EDEF",
X"EFE3",
X"EA84",
X"E98A",
X"EA07",
X"F254",
X"EEE9",
X"F15A",
X"F5BF",
X"F7B3",
X"F6B9",
X"F060",
X"F1D7",
X"FF06",
X"F4C5",
X"FC95",
X"FD12",
X"FAA1",
X"04E2",
X"FD8F",
X"02EE",
X"01F4",
X"05DC",
X"055F",
X"055F",
X"0C35",
X"0B3B",
X"109A",
X"0E29",
X"1117",
X"1405",
X"18E7",
X"1CCF",
X"157C",
X"1FBD",
X"16F3",
X"249F",
X"251C",
X"1A5E",
X"2E63",
X"249F",
X"2616",
X"2693",
X"2BF2",
X"2E63",
X"2BF2",
X"2616",
X"2CEC",
X"2BF2",
X"2887",
X"2D69",
X"2A7B",
X"278D",
X"2D69",
X"249F",
X"2AF8",
X"23A5",
X"251C",
X"2328",
X"15F9",
X"2134",
X"1964",
X"19E1",
X"130B",
X"0F23",
X"0C35",
X"04E2",
X"0177",
X"FE0C",
X"FE0C",
X"FA24",
X"F2D1",
X"F254",
X"EB7E",
X"EEE9",
X"EBFB",
X"F060",
X"F2D1",
X"EB7E",
X"EF66",
X"E90D",
X"EB7E",
X"EA07",
X"E719",
X"E719",
X"E4A8",
X"E525",
X"E890",
X"E890",
X"DE4F",
X"DD55",
X"E61F",
X"DECC",
X"E61F",
X"E890",
X"FA24",
X"EDEF",
X"F3CB",
X"F4C5",
X"EFE3",
X"EA84",
X"E69C",
X"EE6C",
X"EC78",
X"ED72",
X"F254",
X"F4C5",
X"F542",
X"F448",
X"F4C5",
X"FB9B",
X"F34E",
X"F8AD",
X"FC95",
X"0000",
X"FE89",
X"036B",
X"09C4",
X"1194",
X"06D6",
X"0659",
X"05DC",
X"0A41",
X"01F4",
X"0659",
X"0FA0",
X"08CA",
X"0947",
X"03E8",
X"0A41",
X"0271",
X"FD8F",
X"0A41",
X"0659",
X"0753",
X"0465",
X"0CB2",
X"055F",
X"0177",
X"0FA0",
X"08CA",
X"0BB8",
X"0FA0",
X"084D",
X"084D",
X"1194",
X"0DAC",
X"1405",
X"06D6",
X"0ABE",
X"17ED",
X"1194",
X"084D",
X"0659",
X"01F4",
X"F63C",
X"F8AD",
X"ED72",
X"EB01",
X"ED72",
X"E525",
X"E719",
X"E3AE",
X"E4A8",
X"E98A",
X"E90D",
X"E890",
X"E69C",
X"E69C",
X"ED72",
X"EDEF",
X"F3CB",
X"F34E",
X"F7B3",
X"F3CB",
X"F4C5",
X"FF83",
X"FF83",
X"FF83",
X"02EE",
X"07D0",
X"02EE",
X"036B",
X"0659",
X"FE89",
X"FD12",
X"055F",
X"00FA",
X"0659",
X"0753",
X"08CA",
X"0E29",
X"130B",
X"1482",
X"1388",
X"0ABE",
X"0E29",
X"1194",
X"FC18",
X"084D",
X"FF06",
X"FC18",
X"08CA",
X"F830",
X"FF83",
X"0D2F",
X"0947",
X"06D6",
X"0753",
X"0BB8",
X"0E29",
X"1482",
X"0FA0",
X"0D2F",
X"0CB2",
X"0BB8",
X"1211",
X"084D",
X"0ABE",
X"0C35",
X"0271",
X"02EE",
X"02EE",
X"00FA",
X"0D2F",
X"FC95",
X"F6B9",
X"F2D1",
X"E98A",
X"EA07",
X"E525",
X"E3AE",
X"DFC6",
X"DDD2",
X"EA84",
X"E3AE",
X"DAE4",
X"E4A8",
X"D9EA",
X"E2B4",
X"DF49",
X"D8F0",
X"DA67",
X"CF2C",
X"DD55",
X"D67F",
X"DECC",
X"D602",
X"DDD2",
X"DF49",
X"D585",
X"DFC6",
X"DBDE",
X"DBDE",
X"D9EA",
X"E1BA",
X"E13D",
X"DF49",
X"D6FC",
X"DBDE",
X"DA67",
X"D19D",
X"E13D",
X"DAE4",
X"D297",
X"DC5B",
X"DCD8",
X"DDD2",
X"EC78",
X"E61F",
X"DDD2",
X"E525",
X"EBFB",
X"EB7E",
X"EBFB",
X"EB01",
X"EE6C",
X"EBFB",
X"F060",
X"FB9B",
X"F0DD",
X"F542",
X"F830",
X"FD12",
X"FF83",
X"02EE",
X"1211",
X"06D6",
X"0FA0",
X"1770",
X"1A5E",
X"19E1",
X"23A5",
X"20B7",
X"278D",
X"278D",
X"2C6F",
X"2C6F",
X"2BF2",
X"2AF8",
X"22AB",
X"2D69",
X"2981",
X"2328",
X"1FBD",
X"2616",
X"2A7B",
X"20B7",
X"280A",
X"280A",
X"2C6F",
X"2A7B",
X"203A",
X"2D69",
X"249F",
X"2134",
X"2599",
X"2693",
X"2981",
X"2C6F",
X"280A",
X"1FBD",
X"1964",
X"1A5E",
X"1964",
X"101D",
X"157C",
X"101D",
X"109A",
X"1482",
X"18E7",
X"15F9",
X"2422",
X"14FF",
X"101D",
X"18E7",
X"08CA",
X"0EA6",
X"0ABE",
X"0B3B",
X"0177",
X"FF06",
X"03E8",
X"FC18",
X"FAA1",
X"FD12",
X"01F4",
X"0465",
X"0000",
X"0DAC",
X"03E8",
X"FB9B",
X"02EE",
X"03E8",
X"0177",
X"FC95",
X"FD12",
X"07D0",
X"FE0C",
X"F34E",
X"E69C",
X"EEE9",
X"E98A",
X"E237",
X"E331",
X"E2B4",
X"E796",
X"DFC6",
X"E3AE",
X"EB7E",
X"EA07",
X"EBFB",
X"EB01",
X"ECF5",
X"E890",
X"EDEF",
X"F1D7",
X"F7B3",
X"F0DD",
X"EDEF",
X"F92A",
X"F3CB",
X"F0DD",
X"E69C",
X"E42B",
X"DCD8",
X"E3AE",
X"E331",
X"E525",
X"F2D1",
X"E525",
X"E61F",
X"EEE9",
X"E813",
X"F34E",
X"EF66",
X"ED72",
X"F830",
X"F542",
X"F34E",
X"F63C",
X"EFE3",
X"F0DD",
X"EEE9",
X"EFE3",
X"E61F",
X"F2D1",
X"F7B3",
X"F2D1",
X"F830",
X"EFE3",
X"F34E",
X"F4C5",
X"F15A",
X"F34E",
X"F15A",
X"F34E",
X"F1D7",
X"F3CB",
X"F6B9",
X"F9A7",
X"F542",
X"F448",
X"F3CB",
X"F34E",
X"FD8F",
X"F4C5",
X"FF06",
X"F830",
X"F5BF",
X"0659",
X"FB1E",
X"FF06",
X"036B",
X"02EE",
X"08CA",
X"0947",
X"02EE",
X"05DC",
X"FF06",
X"FB9B",
X"05DC",
X"00FA",
X"FE0C",
X"0BB8",
X"0BB8",
X"08CA",
X"1211",
X"1482",
X"128E",
X"109A",
X"16F3",
X"1676",
X"1388",
X"1676",
X"1EC3",
X"2422",
X"2981",
X"2710",
X"1CCF",
X"31CE",
X"251C",
X"278D",
X"2710",
X"2616",
X"22AB",
X"1CCF",
X"2693",
X"2710",
X"2693",
X"2904",
X"1C52",
X"1A5E",
X"1E46",
X"2422",
X"1BD5",
X"15F9",
X"2616",
X"1ADB",
X"186A",
X"14FF",
X"07D0",
X"1388",
X"0E29",
X"09C4",
X"0F23",
X"06D6",
X"1388",
X"1117",
X"1BD5",
X"0FA0",
X"1194",
X"1194",
X"0947",
X"101D",
X"0177",
X"0DAC",
X"03E8",
X"01F4",
X"0DAC",
X"007D",
X"FAA1",
X"FD8F",
X"F4C5",
X"0177",
X"007D",
X"0B3B",
X"0D2F",
X"0947",
X"20B7",
X"19E1",
X"1964",
X"1BD5",
X"16F3",
X"1F40",
X"19E1",
X"157C",
X"1C52",
X"101D",
X"109A",
X"0ABE",
X"02EE",
X"084D",
X"02EE",
X"0BB8",
X"0BB8",
X"04E2",
X"01F4",
X"01F4",
X"F830",
X"FE89",
X"FC95",
X"F6B9",
X"F8AD",
X"F63C",
X"0465",
X"FB9B",
X"0659",
X"0177",
X"0465",
X"FA24",
X"F8AD",
X"084D",
X"FB9B",
X"FB9B",
X"0177",
X"F8AD",
X"FAA1",
X"F15A",
X"EEE9",
X"F92A",
X"ECF5",
X"EEE9",
X"E98A",
X"EC78",
X"EDEF",
X"F060",
X"EFE3",
X"EB7E",
X"EA84",
X"E3AE",
X"E796",
X"E61F",
X"E890",
X"EFE3",
X"EBFB",
X"F7B3",
X"F5BF",
X"F542",
X"FC95",
X"F63C",
X"FB1E",
X"F736",
X"F34E",
X"F060",
X"ECF5",
X"FB1E",
X"F34E",
X"F2D1",
X"F63C",
X"EDEF",
X"FA24",
X"F1D7",
X"ECF5",
X"F5BF",
X"EF66",
X"F1D7",
X"F448",
X"FC18",
X"0947",
X"04E2",
X"02EE",
X"0947",
X"02EE",
X"02EE",
X"FF06",
X"FE0C",
X"FB1E",
X"F542",
X"F060",
X"F34E",
X"EFE3",
X"EC78",
X"EFE3",
X"F15A",
X"F254",
X"EF66",
X"EEE9",
X"ED72",
X"EF66",
X"F0DD",
X"ED72",
X"F060",
X"EC78",
X"EB7E",
X"ED72",
X"F15A",
X"F1D7",
X"F1D7",
X"F060",
X"ED72",
X"EA07",
X"EFE3",
X"ECF5",
X"EEE9",
X"ED72",
X"EA84",
X"ECF5",
X"E796",
X"E813",
X"E4A8",
X"E331",
X"E2B4",
X"DDD2",
X"DECC",
X"E043",
X"E13D",
X"D96D",
X"D96D",
X"D779",
X"D40E",
X"D0A3",
X"CF2C",
X"D67F",
X"DC5B",
X"DAE4",
X"DFC6",
X"D508",
X"DF49",
X"DCD8",
X"DBDE",
X"DC5B",
X"DA67",
X"DECC",
X"DF49",
X"DF49",
X"E4A8",
X"E2B4",
X"E61F",
X"EE6C",
X"E4A8",
X"E719",
X"F736",
X"F8AD",
X"F92A",
X"F9A7",
X"FF06",
X"036B",
X"036B",
X"0000",
X"09C4",
X"055F",
X"05DC",
X"05DC",
X"06D6",
X"0ABE",
X"0EA6",
X"0ABE",
X"0BB8",
X"08CA",
X"007D",
X"0465",
X"09C4",
X"07D0",
X"08CA",
X"0659",
X"0659",
X"04E2",
X"02EE",
X"FD8F",
X"03E8",
X"0947",
X"FD8F",
X"07D0",
X"0CB2",
X"07D0",
X"0D2F",
X"0F23",
X"1CCF",
X"15F9",
X"1194",
X"1117",
X"1A5E",
X"186A",
X"203A",
X"1C52",
X"2328",
X"1964",
X"1BD5",
X"1FBD",
X"2328",
X"278D",
X"2134",
X"2D69",
X"2599",
X"2AF8",
X"32C8",
X"3633",
X"34BC",
X"2F5D",
X"3539",
X"324B",
X"372D",
X"33C2",
X"30D4",
X"30D4",
X"2599",
X"280A",
X"2710",
X"249F",
X"2EE0",
X"2710",
X"2710",
X"2E63",
X"2616",
X"2981",
X"1D4C",
X"251C",
X"1E46",
X"1EC3",
X"1D4C",
X"1B58",
X"1FBD",
X"1A5E",
X"18E7",
X"19E1",
X"1A5E",
X"2328",
X"1ADB",
X"20B7",
X"186A",
X"1F40",
X"1A5E",
X"1C52",
X"222E",
X"1770",
X"2710",
X"23A5",
X"2CEC",
X"2887",
X"2904",
X"23A5",
X"2CEC",
X"203A",
X"1FBD",
X"21B1",
X"1CCF",
X"22AB",
X"2134",
X"2328",
X"1DC9",
X"1BD5",
X"2710",
X"280A",
X"2422",
X"2693",
X"2BF2",
X"2904",
X"23A5",
X"2134",
X"203A",
X"1964",
X"1E46",
X"186A",
X"186A",
X"1482",
X"128E",
X"1194",
X"084D",
X"0ABE",
X"04E2",
X"0177",
X"FE0C",
X"F3CB",
X"F4C5",
X"F7B3",
X"E90D",
X"EFE3",
X"E4A8",
X"E043",
X"E69C",
X"E237",
X"DFC6",
X"DAE4",
X"DF49",
X"D508",
X"DE4F",
X"D779",
X"DA67",
X"D026",
X"D585",
X"DC5B",
X"CDB5",
X"D602",
X"D21A",
X"CA4A",
X"CD38",
X"C6DF",
X"CAC7",
X"C568",
X"C662",
X"CAC7",
X"C568",
X"CBC1",
X"C9CD",
X"CBC1",
X"D297",
X"C950",
X"D19D",
X"D40E",
X"CBC1",
X"D19D",
X"C950",
X"D026",
X"D391",
X"D314",
X"D40E",
X"D8F0",
X"D40E",
X"DB61",
X"DECC",
X"E4A8",
X"DCD8",
X"DECC",
X"DE4F",
X"E525",
X"E42B",
X"E237",
X"E61F",
X"DCD8",
X"E5A2",
X"ECF5",
X"EA07",
X"EA07",
X"E69C",
X"E0C0",
X"ECF5",
X"E98A",
X"EE6C",
X"F1D7",
X"EA84",
X"EFE3",
X"EBFB",
X"F3CB",
X"EEE9",
X"F9A7",
X"F8AD",
X"EEE9",
X"FF83",
X"EF66",
X"EFE3",
X"FAA1",
X"F060",
X"FD12",
X"F9A7",
X"0271",
X"01F4",
X"FC95",
X"0753",
X"F830",
X"F9A7",
X"01F4",
X"F254",
X"FD12",
X"EFE3",
X"E90D",
X"FB1E",
X"EA84",
X"FB1E",
X"FE0C",
X"FA24",
X"0177",
X"0271",
X"0271",
X"0C35",
X"036B",
X"0B3B",
X"08CA",
X"06D6",
X"0B3B",
X"0177",
X"FD8F",
X"03E8",
X"04E2",
X"036B",
X"08CA",
X"09C4",
X"0C35",
X"1ADB",
X"1ADB",
X"2616",
X"20B7",
X"1B58",
X"251C",
X"2134",
X"249F",
X"2B75",
X"2599",
X"2887",
X"2616",
X"23A5",
X"2CEC",
X"2D69",
X"280A",
X"2BF2",
X"2AF8",
X"2C6F",
X"30D4",
X"2EE0",
X"2FDA",
X"2D69",
X"343F",
X"30D4",
X"36B0",
X"2F5D",
X"2FDA",
X"324B",
X"2CEC",
X"2D69",
X"2A7B",
X"2E63",
X"2A7B",
X"2887",
X"2BF2",
X"251C",
X"186A",
X"1B58",
X"23A5",
X"1C52",
X"20B7",
X"21B1",
X"186A",
X"1A5E",
X"1770",
X"14FF",
X"16F3",
X"1388",
X"1405",
X"09C4",
X"036B",
X"0ABE",
X"07D0",
X"0271",
X"01F4",
X"04E2",
X"FE0C",
X"F9A7",
X"F830",
X"0271",
X"055F",
X"0271",
X"0000",
X"F8AD",
X"F2D1",
X"F15A",
X"F254",
X"F34E",
X"007D",
X"007D",
X"00FA",
X"FA24",
X"F63C",
X"F448",
X"EDEF",
X"F63C",
X"E98A",
X"EB7E",
X"E4A8",
X"E90D",
X"F15A",
X"EC78",
X"F3CB",
X"EEE9",
X"E61F",
X"EBFB",
X"EB01",
X"EA07",
X"EA07",
X"EB7E",
X"EF66",
X"E813",
X"E61F",
X"E42B",
X"E331",
X"EB7E",
X"DC5B",
X"E13D",
X"E525",
X"DC5B",
X"E719",
X"D48B",
X"D508",
X"CE32",
X"D120",
X"D67F",
X"D314",
X"D314",
X"D0A3",
X"D508",
X"D602",
X"DA67",
X"D6FC",
X"D297",
X"CE32",
X"D297",
X"D8F0",
X"D96D",
X"D873",
X"D585",
X"D779",
X"D391",
X"D21A",
X"D602",
X"D585",
X"D120",
X"CF2C",
X"D120",
X"D779",
X"DCD8",
X"E69C",
X"E719",
X"E043",
X"E4A8",
X"EC78",
X"E719",
X"DFC6",
X"E0C0",
X"E5A2",
X"E90D",
X"EA84",
X"F736",
X"FE89",
X"FE89",
X"01F4",
X"FE0C",
X"0000",
X"FAA1",
X"F830",
X"F9A7",
X"FAA1",
X"F830",
X"FB9B",
X"00FA",
X"F1D7",
X"F542",
X"F736",
X"FAA1",
X"F448",
X"F15A",
X"F92A",
X"FB1E",
X"03E8",
X"04E2",
X"FC18",
X"FC18",
X"FF06",
X"FF06",
X"FF06",
X"06D6",
X"06D6",
X"084D",
X"130B",
X"084D",
X"101D",
X"1482",
X"15F9",
X"15F9",
X"15F9",
X"278D",
X"21B1",
X"23A5",
X"2710",
X"2693",
X"1BD5",
X"2616",
X"2693",
X"20B7",
X"1EC3",
X"1ADB",
X"222E",
X"15F9",
X"1964",
X"1676",
X"0947",
X"0D2F",
X"0BB8",
X"0F23",
X"0EA6",
X"128E",
X"0ABE",
X"0753",
X"09C4",
X"0947",
X"0CB2",
X"0B3B",
X"0B3B",
X"084D",
X"084D",
X"130B",
X"1770",
X"1194",
X"1676",
X"0DAC",
X"15F9",
X"1405",
X"1964",
X"1D4C",
X"1BD5",
X"222E",
X"22AB",
X"249F",
X"22AB",
X"2B75",
X"203A",
X"249F",
X"23A5",
X"2422",
X"251C",
X"1D4C",
X"1F40",
X"203A",
X"2134",
X"2134",
X"2616",
X"222E",
X"2693",
X"2693",
X"20B7",
X"1FBD",
X"2693",
X"2328",
X"1C52",
X"2422",
X"186A",
X"0F23",
X"0EA6",
X"09C4",
X"128E",
X"084D",
X"0947",
X"0EA6",
X"0A41",
X"0ABE",
X"109A",
X"055F",
X"05DC",
X"0C35",
X"03E8",
X"055F",
X"09C4",
X"0EA6",
X"1482",
X"0F23",
X"0BB8",
X"0659",
X"09C4",
X"FE89",
X"F736",
X"FD8F",
X"03E8",
X"F63C",
X"FF06",
X"F63C",
X"FA24",
X"F9A7",
X"F3CB",
X"F34E",
X"F448",
X"FB9B",
X"F736",
X"FF83",
X"FA24",
X"F8AD",
X"FD8F",
X"F92A",
X"F7B3",
X"F830",
X"FB1E",
X"F9A7",
X"FC95",
X"FB9B",
X"FC18",
X"0177",
X"FC95",
X"FC95",
X"FF06",
X"F9A7",
X"FB1E",
X"F7B3",
X"F92A",
X"FB1E",
X"F736",
X"F7B3",
X"FC95",
X"0177",
X"FD12",
X"01F4",
X"00FA",
X"084D",
X"FD12",
X"007D",
X"04E2",
X"0271",
X"0C35",
X"00FA",
X"09C4",
X"0753",
X"007D",
X"0271",
X"F6B9",
X"F830",
X"F3CB",
X"F736",
X"F34E",
X"EB01",
X"E69C",
X"E3AE",
X"E2B4",
X"E2B4",
X"DC5B",
X"DCD8",
X"DA67",
X"D48B",
X"D96D",
X"D391",
X"D7F6",
X"D96D",
X"D6FC",
X"DD55",
X"DC5B",
X"DB61",
X"D873",
X"D6FC",
X"D297",
X"D873",
X"DC5B",
X"DFC6",
X"E043",
X"DBDE",
X"E237",
X"DF49",
X"D96D",
X"DAE4",
X"E5A2",
X"DF49",
X"DB61",
X"E3AE",
X"E61F",
X"E5A2",
X"EB01",
X"F5BF",
X"F9A7",
X"F15A",
X"F9A7",
X"036B",
X"FC18",
X"FE0C",
X"0753",
X"0465",
X"0DAC",
X"1405",
X"1770",
X"1D4C",
X"1211",
X"1EC3",
X"1A5E",
X"1CCF",
X"21B1",
X"2887",
X"2981",
X"2F5D",
X"2E63",
X"3345",
X"3539",
X"3345",
X"3151",
X"324B",
X"30D4",
X"29FE",
X"2DE6",
X"30D4",
X"33C2",
X"3345",
X"32C8",
X"35B6",
X"2B75",
X"2A7B",
X"2710",
X"2710",
X"222E",
X"1BD5",
X"1E46",
X"1D4C",
X"1DC9",
X"1BD5",
X"1CCF",
X"17ED",
X"17ED",
X"1676",
X"17ED",
X"18E7",
X"18E7",
X"1B58",
X"16F3",
X"15F9",
X"109A",
X"0A41",
X"0A41",
X"0465",
X"05DC",
X"09C4",
X"00FA",
X"FF83",
X"F830",
X"EE6C",
X"ED72",
X"E813",
X"E42B",
X"E4A8",
X"DDD2",
X"DDD2",
X"DC5B",
X"DDD2",
X"DECC",
X"DAE4",
X"DF49",
X"D40E",
X"D602",
X"D6FC",
X"D0A3",
X"D21A",
X"CDB5",
X"C9CD",
X"C856",
X"C6DF",
X"CBC1",
X"C9CD",
X"C9CD",
X"CC3E",
X"CB44",
X"CDB5",
X"CC3E",
X"D297",
X"D21A",
X"D40E",
X"D120",
X"D21A",
X"D297",
X"DAE4",
X"D602",
X"D779",
X"DAE4",
X"D96D",
X"DC5B",
X"DA67",
X"DDD2",
X"DA67",
X"CFA9",
X"D602",
X"D873",
X"DBDE",
X"DD55",
X"E331",
X"E890",
X"EA84",
X"F2D1",
X"F4C5",
X"F9A7",
X"01F4",
X"0465",
X"FC95",
X"FB9B",
X"FF06",
X"FD8F",
X"036B",
X"06D6",
X"08CA",
X"0CB2",
X"0FA0",
X"157C",
X"128E",
X"19E1",
X"101D",
X"0DAC",
X"0CB2",
X"0CB2",
X"0B3B",
X"0D2F",
X"128E",
X"0659",
X"FF83",
X"02EE",
X"06D6",
X"0947",
X"0465",
X"FD12",
X"0177",
X"00FA",
X"00FA",
X"084D",
X"0B3B",
X"0465",
X"0753",
X"084D",
X"07D0",
X"03E8",
X"FC95",
X"03E8",
X"0000",
X"FF06",
X"01F4",
X"FF06",
X"04E2",
X"FB1E",
X"00FA",
X"04E2",
X"07D0",
X"0947",
X"084D",
X"0C35",
X"06D6",
X"0BB8",
X"0EA6",
X"0D2F",
X"0D2F",
X"128E",
X"0BB8",
X"084D",
X"084D",
X"06D6",
X"08CA",
X"FB9B",
X"0271",
X"FD12",
X"036B",
X"FE0C",
X"F7B3",
X"FE0C",
X"FB9B",
X"FA24",
X"F736",
X"F2D1",
X"F4C5",
X"F7B3",
X"ED72",
X"EBFB",
X"EF66",
X"EF66",
X"007D",
X"FC95",
X"FF83",
X"FB1E",
X"FF06",
X"03E8",
X"04E2",
X"0CB2",
X"07D0",
X"06D6",
X"08CA",
X"07D0",
X"03E8",
X"0B3B",
X"0BB8",
X"0EA6",
X"0C35",
X"0FA0",
X"14FF",
X"0FA0",
X"1117",
X"0E29",
X"1211",
X"1BD5",
X"1CCF",
X"14FF",
X"16F3",
X"1CCF",
X"17ED",
X"1F40",
X"1A5E",
X"1D4C",
X"249F",
X"1BD5",
X"2134",
X"23A5",
X"2599",
X"278D",
X"251C",
X"2599",
X"2EE0",
X"2CEC",
X"2E63",
X"3151",
X"2F5D",
X"2DE6",
X"3057",
X"3057",
X"29FE",
X"3057",
X"2AF8",
X"2BF2",
X"278D",
X"2710",
X"2BF2",
X"2616",
X"2B75",
X"2328",
X"2EE0",
X"222E",
X"2710",
X"2AF8",
X"2328",
X"1F40",
X"1D4C",
X"18E7",
X"14FF",
X"14FF",
X"1388",
X"15F9",
X"0F23",
X"09C4",
X"084D",
X"08CA",
X"036B",
X"084D",
X"01F4",
X"0000",
X"FB9B",
X"F830",
X"FC95",
X"F8AD",
X"F4C5",
X"EC78",
X"EFE3",
X"EB01",
X"EC78",
X"EBFB",
X"E90D",
X"E719",
X"E890",
X"DF49",
X"E90D",
X"E2B4",
X"DFC6",
X"E69C",
X"E813",
X"E61F",
X"E4A8",
X"E98A",
X"E813",
X"ED72",
X"F5BF",
X"F060",
X"F1D7",
X"F3CB",
X"F254",
X"FD8F",
X"F254",
X"F2D1",
X"F63C",
X"F448",
X"EA84",
X"F1D7",
X"F830",
X"F63C",
X"F3CB",
X"F92A",
X"FE89",
X"F254",
X"FB9B",
X"F830",
X"F7B3",
X"F63C",
X"F63C",
X"FB9B",
X"F7B3",
X"F63C",
X"F5BF",
X"F34E",
X"FA24",
X"F92A",
X"F542",
X"F736",
X"F7B3",
X"F6B9",
X"F830",
X"F7B3",
X"F9A7",
X"FB1E",
X"FAA1",
X"FB9B",
X"F542",
X"FAA1",
X"FB1E",
X"F9A7",
X"FC18",
X"F63C",
X"FE0C",
X"FC18",
X"FB9B",
X"FC95",
X"FC95",
X"FA24",
X"F0DD",
X"FD12",
X"F34E",
X"F0DD",
X"F736",
X"FA24",
X"F34E",
X"F4C5",
X"F7B3",
X"FF83",
X"F92A",
X"F3CB",
X"ECF5",
X"E719",
X"F15A",
X"E3AE",
X"EB7E",
X"E525",
X"E1BA",
X"E043",
X"E237",
X"E719",
X"E42B",
X"E13D",
X"E3AE",
X"E13D",
X"E796",
X"E525",
X"E890",
X"ED72",
X"E813",
X"E890",
X"E90D",
X"E796",
X"E813",
X"EB7E",
X"E890",
X"EB7E",
X"EDEF",
X"EC78",
X"ED72",
X"F0DD",
X"F254",
X"F5BF",
X"F3CB",
X"EFE3",
X"F1D7",
X"F254",
X"F5BF",
X"F736",
X"F5BF",
X"F7B3",
X"EF66",
X"F448",
X"F6B9",
X"F63C",
X"F6B9",
X"F254",
X"F92A",
X"F7B3",
X"F5BF",
X"FB1E",
X"03E8",
X"03E8",
X"0659",
X"084D",
X"04E2",
X"03E8",
X"00FA",
X"0271",
X"03E8",
X"05DC",
X"04E2",
X"0465",
X"0ABE",
X"04E2",
X"0947",
X"0CB2",
X"09C4",
X"08CA",
X"0DAC",
X"0CB2",
X"0EA6",
X"0EA6",
X"0CB2",
X"0FA0",
X"14FF",
X"1211",
X"1117",
X"0EA6",
X"0FA0",
X"0FA0",
X"1388",
X"130B",
X"109A",
X"1482",
X"1676",
X"1676",
X"1676",
X"18E7",
X"16F3",
X"19E1",
X"1B58",
X"186A",
X"16F3",
X"1482",
X"0FA0",
X"1482",
X"0DAC",
X"109A",
X"0CB2",
X"0C35",
X"07D0",
X"06D6",
X"03E8",
X"0753",
X"FD12",
X"036B",
X"0465",
X"FB1E",
X"01F4",
X"FF83",
X"055F",
X"05DC",
X"02EE",
X"0177",
X"07D0",
X"0659",
X"0271",
X"09C4",
X"0E29",
X"07D0",
X"0E29",
X"0947",
X"07D0",
X"0B3B",
X"07D0",
X"07D0",
X"06D6",
X"0659",
X"0659",
X"06D6",
X"04E2",
X"0659",
X"FE0C",
X"0000",
X"FF83",
X"FAA1",
X"F63C",
X"F3CB",
X"F448",
X"F4C5",
X"EEE9",
X"F34E",
X"EF66",
X"ED72",
X"EB01",
X"EEE9",
X"F0DD",
X"EFE3",
X"F542",
X"F34E",
X"EBFB",
X"F736",
X"F542",
X"F34E",
X"F9A7",
X"F830",
X"F2D1",
X"E98A",
X"EFE3",
X"EF66",
X"F3CB",
X"F1D7",
X"F542",
X"F34E",
X"F8AD",
X"F7B3",
X"F9A7",
X"FF06",
X"FE0C",
X"03E8",
X"F830",
X"007D",
X"F254",
X"F92A",
X"F4C5",
X"E98A",
X"ED72",
X"E42B",
X"E61F",
X"EA07",
X"DB61",
X"E0C0",
X"E043",
X"DDD2",
X"DE4F",
X"D9EA",
X"DECC",
X"E043",
X"E69C",
X"E4A8",
X"E3AE",
X"E796",
X"EEE9",
X"F3CB",
X"F6B9",
X"FB9B",
X"FE89",
X"FAA1",
X"0000",
X"0A41",
X"007D",
X"0BB8",
X"0753",
X"07D0",
X"128E",
X"08CA",
X"186A",
X"0E29",
X"157C",
X"1964",
X"1211",
X"1CCF",
X"186A",
X"1964",
X"1117",
X"0FA0",
X"15F9",
X"0BB8",
X"0B3B",
X"101D",
X"19E1",
X"1FBD",
X"1EC3",
X"1ADB",
X"1E46",
X"1D4C",
X"18E7",
X"249F",
X"1B58",
X"1DC9",
X"1F40",
X"1482",
X"251C",
X"1A5E",
X"2134",
X"23A5",
X"1770",
X"1676",
X"1E46",
X"1770",
X"1194",
X"1482",
X"0C35",
X"157C",
X"0B3B",
X"101D",
X"0B3B",
X"0DAC",
X"0947",
X"084D",
X"04E2",
X"0753",
X"0271",
X"F448",
X"04E2",
X"F9A7",
X"F9A7",
X"FD12",
X"F5BF",
X"F542",
X"F1D7",
X"EF66",
X"F63C",
X"F0DD",
X"E719",
X"ECF5",
X"EA07",
X"EA84",
X"E98A",
X"E98A",
X"EBFB",
X"EBFB",
X"E813",
X"EB01",
X"EEE9",
X"F63C",
X"F63C",
X"F2D1",
X"F9A7",
X"F9A7",
X"FC95",
X"036B",
X"05DC",
X"0177",
X"0465",
X"07D0",
X"0CB2",
X"101D",
X"0CB2",
X"109A",
X"0FA0",
X"130B",
X"1194",
X"1D4C",
X"1964",
X"14FF",
X"157C",
X"101D",
X"14FF",
X"16F3",
X"14FF",
X"17ED",
X"1C52",
X"17ED",
X"19E1",
X"1B58",
X"19E1",
X"1A5E",
X"17ED",
X"157C",
X"0FA0",
X"128E",
X"128E",
X"0F23",
X"128E",
X"14FF",
X"1405",
X"157C",
X"1194",
X"101D",
X"0F23",
X"0E29",
X"0C35",
X"084D",
X"07D0",
X"05DC",
X"07D0",
X"0C35",
X"0659",
X"0ABE",
X"0BB8",
X"0271",
X"02EE",
X"FD12",
X"007D",
X"FC18",
X"FA24",
X"FC95",
X"FE89",
X"FE89",
X"0177",
X"F92A",
X"FC18",
X"F830",
X"F4C5",
X"F6B9",
X"F63C",
X"F6B9",
X"F736",
X"F92A",
X"FC18",
X"FAA1",
X"FB1E",
X"FD12",
X"F448",
X"F830",
X"F8AD",
X"F542",
X"F7B3",
X"FC95",
X"FC95",
X"F9A7",
X"FB9B",
X"FE0C",
X"FD8F",
X"FAA1",
X"FE89",
X"F8AD",
X"F1D7",
X"F736",
X"F8AD",
X"F2D1",
X"F254",
X"EE6C",
X"EEE9",
X"EFE3",
X"ECF5",
X"ED72",
X"EBFB",
X"E796",
X"E813",
X"ECF5",
X"EBFB",
X"EB7E",
X"EFE3",
X"F254",
X"F34E",
X"F5BF",
X"F1D7",
X"F34E",
X"F34E",
X"F1D7",
X"F830",
X"F15A",
X"F34E",
X"F542",
X"EF66",
X"F448",
X"F542",
X"FC95",
X"FB9B",
X"F736",
X"F448",
X"F34E",
X"EDEF",
X"F7B3",
X"F736",
X"F254",
X"F736",
X"F448",
X"007D",
X"FA24",
X"FE0C",
X"FF83",
X"FE0C",
X"FD12",
X"FD12",
X"00FA",
X"0465",
X"03E8",
X"09C4",
X"084D",
X"03E8",
X"08CA",
X"02EE",
X"0A41",
X"0753",
X"01F4",
X"0A41",
X"1194",
X"0B3B",
X"0ABE",
X"1211",
X"0F23",
X"0D2F",
X"0D2F",
X"0F23",
X"0753",
X"0947",
X"15F9",
X"0E29",
X"109A",
X"1117",
X"0CB2",
X"1388",
X"0FA0",
X"128E",
X"109A",
X"101D",
X"0EA6",
X"0659",
X"06D6",
X"084D",
X"0000",
X"09C4",
X"FB1E",
X"055F",
X"02EE",
X"0000",
X"0659",
X"03E8",
X"04E2",
X"04E2",
X"0753",
X"09C4",
X"0659",
X"084D",
X"0271",
X"0659",
X"0753",
X"0000",
X"0947",
X"00FA",
X"FE89",
X"FC95",
X"FB1E",
X"FE0C",
X"FB9B",
X"FC18",
X"F9A7",
X"F7B3",
X"F9A7",
X"FAA1",
X"F4C5",
X"F448",
X"F448",
X"F5BF",
X"F736",
X"F7B3",
X"F34E",
X"F34E",
X"F2D1",
X"F34E",
X"F34E",
X"ECF5",
X"EF66",
X"F34E",
X"EFE3",
X"EA07",
X"E890",
X"E98A",
X"EC78",
X"ECF5",
X"E813",
X"E69C",
X"E331",
X"E813",
X"E3AE",
X"D96D",
X"E1BA",
X"DBDE",
X"D779",
X"D314",
X"D585",
X"D297",
X"D314",
X"D8F0",
X"D40E",
X"CBC1",
X"DCD8",
X"D508",
X"CDB5",
X"D0A3",
X"D19D",
X"D120",
X"D9EA",
X"D19D",
X"D7F6",
X"E043",
X"D9EA",
X"D8F0",
X"DB61",
X"D779",
X"D6FC",
X"D6FC",
X"D779",
X"DAE4",
X"DA67",
X"DBDE",
X"CFA9",
X"DDD2",
X"DE4F",
X"DE4F",
X"E331",
X"E043",
X"E5A2",
X"EE6C",
X"E2B4",
X"E69C",
X"F1D7",
X"EA84",
X"EF66",
X"F63C",
X"EDEF",
X"F2D1",
X"F542",
X"F92A",
X"FA24",
X"007D",
X"FF06",
X"0271",
X"0947",
X"09C4",
X"09C4",
X"0EA6",
X"06D6",
X"0E29",
X"14FF",
X"07D0",
X"0B3B",
X"101D",
X"0C35",
X"1676",
X"157C",
X"157C",
X"1C52",
X"1BD5",
X"1A5E",
X"1964",
X"1A5E",
X"19E1",
X"1DC9",
X"1DC9",
X"19E1",
X"1964",
X"19E1",
X"18E7",
X"1CCF",
X"1A5E",
X"1A5E",
X"1FBD",
X"1C52",
X"1BD5",
X"1CCF",
X"249F",
X"1E46",
X"1C52",
X"1A5E",
X"15F9",
X"1D4C",
X"1211",
X"1676",
X"186A",
X"186A",
X"1964",
X"1964",
X"20B7",
X"1FBD",
X"2422",
X"1FBD",
X"1BD5",
X"2599",
X"2710",
X"278D",
X"2693",
X"2693",
X"2904",
X"278D",
X"2981",
X"2B75",
X"2710",
X"2DE6",
X"2E63",
X"2DE6",
X"3057",
X"30D4",
X"3345",
X"343F",
X"2A7B",
X"2A7B",
X"35B6",
X"2B75",
X"2A7B",
X"35B6",
X"3057",
X"2A7B",
X"2DE6",
X"2DE6",
X"2CEC",
X"2DE6",
X"2AF8",
X"3151",
X"2F5D",
X"2CEC",
X"2DE6",
X"2EE0",
X"2C6F",
X"2AF8",
X"2FDA",
X"2C6F",
X"2CEC",
X"2AF8",
X"2887",
X"280A",
X"278D",
X"2710",
X"278D",
X"2616",
X"280A",
X"2710",
X"1FBD",
X"2693",
X"2599",
X"20B7",
X"249F",
X"1F40",
X"23A5",
X"23A5",
X"1E46",
X"2599",
X"1D4C",
X"1405",
X"1964",
X"1405",
X"109A",
X"0A41",
X"02EE",
X"03E8",
X"036B",
X"07D0",
X"FE89",
X"FA24",
X"F830",
X"F4C5",
X"F254",
X"EC78",
X"F8AD",
X"F254",
X"ED72",
X"E90D",
X"EA84",
X"EB7E",
X"E5A2",
X"E796",
X"E525",
X"E043",
X"DE4F",
X"DC5B",
X"DA67",
X"D779",
X"D508",
X"D6FC",
X"D48B",
X"D508",
X"D585",
X"D21A",
X"D48B",
X"D391",
X"D391",
X"D391",
X"D48B",
X"D7F6",
X"D602",
X"D19D",
X"D19D",
X"D314",
X"D21A",
X"D026",
X"D0A3",
X"D585",
X"CE32",
X"CE32",
X"CE32",
X"CB44",
X"CAC7",
X"CB44",
X"CF2C",
X"C950",
X"C950",
X"CC3E",
X"C8D3",
X"C950",
X"CF2C",
X"D0A3",
X"D297",
X"D026",
X"CD38",
X"C950",
X"D026",
X"CFA9",
X"CBC1",
X"CC3E",
X"D21A",
X"D391",
X"D297",
X"D026",
X"D40E",
X"D67F",
X"D8F0",
X"D7F6",
X"D19D",
X"DAE4",
X"DA67",
X"DBDE",
X"E0C0",
X"E331",
X"E0C0",
X"E2B4",
X"E69C",
X"EA84",
X"EA84",
X"EC78",
X"EDEF",
X"EF66",
X"EEE9",
X"EEE9",
X"F92A",
X"FA24",
X"F736",
X"F7B3",
X"F9A7",
X"F92A",
X"F736",
X"F34E",
X"F6B9",
X"F5BF",
X"F3CB",
X"F3CB",
X"F5BF",
X"F7B3",
X"F736",
X"FC95",
X"FE0C",
X"01F4",
X"0947",
X"0D2F",
X"1388",
X"128E",
X"0D2F",
X"1405",
X"14FF",
X"1388",
X"16F3",
X"1482",
X"1676",
X"1770",
X"157C",
X"1964",
X"1EC3",
X"1A5E",
X"1D4C",
X"20B7",
X"1B58",
X"1B58",
X"1D4C",
X"1D4C",
X"1C52",
X"1F40",
X"222E",
X"1CCF",
X"1D4C",
X"1EC3",
X"1D4C",
X"2422",
X"23A5",
X"2710",
X"2A7B",
X"2981",
X"2A7B",
X"2981",
X"29FE",
X"2981",
X"280A",
X"2E63",
X"2D69",
X"2981",
X"2710",
X"2328",
X"2328",
X"2422",
X"1FBD",
X"1C52",
X"1DC9",
X"1ADB",
X"15F9",
X"14FF",
X"1388",
X"0DAC",
X"0F23",
X"0BB8",
X"08CA",
X"1117",
X"07D0",
X"04E2",
X"055F",
X"00FA",
X"01F4",
X"04E2",
X"FF06",
X"FB9B",
X"FF06",
X"FE0C",
X"FB9B",
X"F92A",
X"F92A",
X"F92A",
X"F7B3",
X"F736",
X"F830",
X"F6B9",
X"F6B9",
X"F4C5",
X"F2D1",
X"F4C5",
X"F6B9",
X"F060",
X"EC78",
X"EB7E",
X"E90D",
X"EA07",
X"E719",
X"E4A8",
X"E525",
X"E525",
X"E0C0",
X"E4A8",
X"E2B4",
X"D9EA",
X"DA67",
X"DBDE",
X"D585",
X"D873",
X"D7F6",
X"D314",
X"D391",
X"D391",
X"D40E",
X"D602",
X"D48B",
X"D19D",
X"D297",
X"D026",
X"D120",
X"D026",
X"CDB5",
X"CDB5",
X"CF2C",
X"D21A",
X"D0A3",
X"CF2C",
X"D67F",
X"D873",
X"D9EA",
X"DC5B",
X"DAE4",
X"DC5B",
X"DFC6",
X"E719",
X"E813",
X"EB01",
X"E98A",
X"ED72",
X"F830",
X"F2D1",
X"F542",
X"FD12",
X"FB1E",
X"0000",
X"07D0",
X"0465",
X"05DC",
X"0FA0",
X"1405",
X"109A",
X"1676",
X"1194",
X"0C35",
X"1676",
X"1388",
X"1482",
X"1B58",
X"1A5E",
X"19E1",
X"1C52",
X"1B58",
X"15F9",
X"157C",
X"17ED",
X"18E7",
X"14FF",
X"19E1",
X"1B58",
X"157C",
X"1C52",
X"1BD5",
X"222E",
X"2422",
X"2710",
X"251C",
X"2422",
X"2693",
X"2887",
X"2E63",
X"2FDA",
X"2FDA",
X"30D4",
X"31CE",
X"3345",
X"33C2",
X"2FDA",
X"2CEC",
X"2A7B",
X"2CEC",
X"3151",
X"2DE6",
X"343F",
X"2B75",
X"3151",
X"3539",
X"2AF8",
X"2AF8",
X"2CEC",
X"2904",
X"2904",
X"2887",
X"2B75",
X"2A7B",
X"2BF2",
X"2EE0",
X"3151",
X"30D4",
X"30D4",
X"2D69",
X"2DE6",
X"2FDA",
X"2B75",
X"2AF8",
X"29FE",
X"2CEC",
X"2C6F",
X"280A",
X"2887",
X"2D69",
X"2A7B",
X"2904",
X"2693",
X"22AB",
X"222E",
X"2422",
X"21B1",
X"222E",
X"2134",
X"21B1",
X"23A5",
X"1DC9",
X"23A5",
X"2134",
X"1F40",
X"1A5E",
X"1770",
X"18E7",
X"16F3",
X"16F3",
X"1676",
X"1482",
X"1676",
X"130B",
X"1405",
X"1770",
X"1211",
X"1194",
X"101D",
X"1194",
X"1770",
X"109A",
X"128E",
X"1405",
X"0FA0",
X"0CB2",
X"0A41",
X"02EE",
X"01F4",
X"0000",
X"F6B9",
X"F63C",
X"F92A",
X"ED72",
X"F7B3",
X"F2D1",
X"EA84",
X"EF66",
X"EB01",
X"EB01",
X"E4A8",
X"E719",
X"E61F",
X"DCD8",
X"DAE4",
X"E13D",
X"E1BA",
X"E42B",
X"E043",
X"DBDE",
X"DDD2",
X"D9EA",
X"D9EA",
X"D67F",
X"D585",
X"D120",
X"CEAF",
X"CA4A",
X"D026",
X"D21A",
X"D0A3",
X"D391",
X"D602",
X"CE32",
X"D19D",
X"D602",
X"C8D3",
X"D19D",
X"C6DF",
X"CC3E",
X"D026",
X"C9CD",
X"D026",
X"CF2C",
X"D391",
X"CF2C",
X"D19D",
X"D026",
X"CDB5",
X"CD38",
X"CAC7",
X"CFA9",
X"CDB5",
X"D026",
X"D297",
X"CB44",
X"CEAF",
X"CD38",
X"CBC1",
X"D391",
X"CE32",
X"C9CD",
X"CBC1",
X"CD38",
X"CBC1",
X"CAC7",
X"CE32",
X"D026",
X"CFA9",
X"D026",
X"D0A3",
X"D0A3",
X"D67F",
X"D297",
X"D19D",
X"D19D",
X"D508",
X"D6FC",
X"D6FC",
X"D9EA",
X"DD55",
X"E0C0",
X"DD55",
X"DECC",
X"E42B",
X"E61F",
X"E42B",
X"E813",
X"EA84",
X"EA84",
X"EB01",
X"EEE9",
X"F5BF",
X"F7B3",
X"FB1E",
X"FC18",
X"01F4",
X"03E8",
X"0753",
X"0947",
X"0753",
X"0CB2",
X"0F23",
X"101D",
X"157C",
X"1388",
X"157C",
X"1482",
X"1676",
X"1482",
X"128E",
X"0F23",
X"0BB8",
X"0CB2",
X"084D",
X"07D0",
X"0B3B",
X"08CA",
X"09C4",
X"08CA",
X"0A41",
X"0BB8",
X"0ABE",
X"0B3B",
X"06D6",
X"0DAC",
X"0C35",
X"0ABE",
X"09C4",
X"0EA6",
X"109A",
X"1117",
X"1211",
X"1194",
X"0F23",
X"130B",
X"1405",
X"0FA0",
X"1194",
X"1770",
X"17ED",
X"1770",
X"1E46",
X"23A5",
X"2710",
X"2981",
X"2B75",
X"2DE6",
X"2DE6",
X"2E63",
X"2F5D",
X"2F5D",
X"2E63",
X"31CE",
X"2FDA",
X"2DE6",
X"2BF2",
X"2DE6",
X"2EE0",
X"2DE6",
X"2C6F",
X"2EE0",
X"324B",
X"35B6",
X"31CE",
X"324B",
X"2F5D",
X"2AF8",
X"2B75",
X"3057",
X"31CE",
X"30D4",
X"2EE0",
X"2DE6",
X"3151",
X"33C2",
X"30D4",
X"2F5D",
X"2C6F",
X"2CEC",
X"2DE6",
X"2BF2",
X"2B75",
X"2CEC",
X"2AF8",
X"2E63",
X"2D69",
X"2887",
X"2981",
X"251C",
X"2616",
X"21B1",
X"2693",
X"249F",
X"1DC9",
X"1FBD",
X"1964",
X"17ED",
X"157C",
X"1211",
X"14FF",
X"128E",
X"0A41",
X"0B3B",
X"0ABE",
X"06D6",
X"03E8",
X"02EE",
X"FC18",
X"F9A7",
X"F6B9",
X"F448",
X"F736",
X"EDEF",
X"E61F",
X"E42B",
X"DDD2",
X"D96D",
X"D96D",
X"D0A3",
X"D585",
X"D6FC",
X"D391",
X"CDB5",
X"CA4A",
X"CC3E",
X"C950",
X"C5E5",
X"CBC1",
X"C4EB",
X"C5E5",
X"C8D3",
X"C5E5",
X"C8D3",
X"C5E5",
X"C6DF",
X"C8D3",
X"C5E5",
X"C9CD",
X"CBC1",
X"CB44",
X"CCBB",
X"C856",
X"C75C",
X"CC3E",
X"CBC1",
X"CD38",
X"D0A3",
X"D297",
X"CAC7",
X"CB44",
X"D026",
X"CE32",
X"CEAF",
X"D120",
X"CE32",
X"D0A3",
X"D314",
X"D602",
X"D508",
X"D96D",
X"DB61",
X"D7F6",
X"D67F",
X"D6FC",
X"D7F6",
X"D8F0",
X"D96D",
X"DB61",
X"DC5B",
X"DAE4",
X"DECC",
X"E0C0",
X"DFC6",
X"DECC",
X"DCD8",
X"DE4F",
X"E043",
X"E1BA",
X"E3AE",
X"E42B",
X"E525",
X"E813",
X"E69C",
X"EA07",
X"EA84",
X"EB01",
X"EBFB",
X"E90D",
X"EC78",
X"EE6C",
X"F15A",
X"F2D1",
X"F448",
X"F34E",
X"EEE9",
X"F1D7",
X"F34E",
X"F060",
X"F15A",
X"F2D1",
X"F3CB",
X"F4C5",
X"F736",
X"F5BF",
X"F5BF",
X"FAA1",
X"F92A",
X"F63C",
X"F92A",
X"FE89",
X"FE89",
X"FD8F",
X"0177",
X"007D",
X"0465",
X"055F",
X"0A41",
X"101D",
X"15F9",
X"157C",
X"17ED",
X"1BD5",
X"222E",
X"2422",
X"278D",
X"2887",
X"2AF8",
X"2FDA",
X"2FDA",
X"324B",
X"36B0",
X"372D",
X"3827",
X"34BC",
X"3633",
X"38A4",
X"3539",
X"343F",
X"35B6",
X"3539",
X"37AA",
X"372D",
X"38A4",
X"3B15",
X"37AA",
X"3B15",
X"37AA",
X"3633",
X"343F",
X"37AA",
X"3539",
X"3539",
X"35B6",
X"33C2",
X"324B",
X"36B0",
X"3633",
X"2F5D",
X"343F",
X"372D",
X"33C2",
X"32C8",
X"3151",
X"324B",
X"30D4",
X"2EE0",
X"2FDA",
X"2E63",
X"2CEC",
X"2B75",
X"2BF2",
X"280A",
X"2C6F",
X"2BF2",
X"2599",
X"2422",
X"20B7",
X"2616",
X"1D4C",
X"1A5E",
X"1DC9",
X"1BD5",
X"1ADB",
X"1A5E",
X"1E46",
X"16F3",
X"14FF",
X"0E29",
X"1117",
X"0EA6",
X"0DAC",
X"0A41",
X"055F",
X"03E8",
X"0000",
X"007D",
X"FAA1",
X"FB1E",
X"FF83",
X"F830",
X"F6B9",
X"F254",
X"F34E",
X"F3CB",
X"E890",
X"E796",
X"EE6C",
X"EA07",
X"E813",
X"E61F",
X"E1BA",
X"E890",
X"E331",
X"E4A8",
X"E42B",
X"DB61",
X"E043",
X"DF49",
X"DB61",
X"D96D",
X"D8F0",
X"D602",
X"D67F",
X"D297",
X"D602",
X"D314",
X"D314",
X"D508",
X"D120",
X"D40E",
X"D508",
X"CF2C",
X"CDB5",
X"D779",
X"D508",
X"D19D",
X"D508",
X"CCBB",
X"CDB5",
X"D0A3",
X"D314",
X"D40E",
X"D120",
X"D508",
X"D508",
X"D67F",
X"D873",
X"DBDE",
X"D8F0",
X"D602",
X"D0A3",
X"D585",
X"D120",
X"D48B",
X"D585",
X"D297",
X"D508",
X"CCBB",
X"D19D",
X"D19D",
X"D314",
X"D21A",
X"D120",
X"D21A",
X"D21A",
X"D120",
X"D391",
X"D602",
X"D67F",
X"D602",
X"DC5B",
X"DA67",
X"DA67",
X"E043",
X"DE4F",
X"E1BA",
X"E043",
X"E13D",
X"E4A8",
X"DE4F",
X"E0C0",
X"E2B4",
X"E13D",
X"E237",
X"DECC",
X"E1BA",
X"E1BA",
X"E043",
X"EBFB",
X"E331",
X"E796",
X"E719",
X"E4A8",
X"DFC6",
X"E719",
X"E525",
X"E69C",
X"ECF5",
X"EA84",
X"F254",
X"EDEF",
X"EDEF",
X"EDEF",
X"F3CB",
X"F448",
X"EE6C",
X"ED72",
X"F63C",
X"F060",
X"F3CB",
X"F736",
X"FC95",
X"0000",
X"F830",
X"FE0C",
X"07D0",
X"0FA0",
X"1117",
X"1964",
X"186A",
X"1E46",
X"1DC9",
X"1FBD",
X"2A7B",
X"2710",
X"2981",
X"2B75",
X"2710",
X"2693",
X"2887",
X"2C6F",
X"2EE0",
X"2AF8",
X"32C8",
X"3827",
X"35B6",
X"33C2",
X"3A1B",
X"3B92",
X"372D",
X"3921",
X"3827",
X"343F",
X"3921",
X"3A98",
X"36B0",
X"3539",
X"37AA",
X"399E",
X"372D",
X"399E",
X"343F",
X"3921",
X"3151",
X"324B",
X"372D",
X"2EE0",
X"38A4",
X"372D",
X"3057",
X"2CEC",
X"2F5D",
X"2FDA",
X"2EE0",
X"2EE0",
X"2DE6",
X"2BF2",
X"2BF2",
X"324B",
X"2F5D",
X"2B75",
X"2B75",
X"2904",
X"2887",
X"2693",
X"22AB",
X"249F",
X"251C",
X"2599",
X"222E",
X"1C52",
X"1EC3",
X"2134",
X"1D4C",
X"1482",
X"1964",
X"130B",
X"109A",
X"0C35",
X"0C35",
X"0753",
X"00FA",
X"0465",
X"06D6",
X"0465",
X"00FA",
X"00FA",
X"FD8F",
X"FD12",
X"FD12",
X"F448",
X"F448",
X"F4C5",
X"EE6C",
X"EDEF",
X"EA07",
X"E90D",
X"E331",
X"E1BA",
X"DCD8",
X"D96D",
X"DDD2",
X"DE4F",
X"E525",
X"E1BA",
X"E4A8",
X"EA07",
X"EDEF",
X"F2D1",
X"F92A",
X"F9A7",
X"F92A",
X"FD8F",
X"036B",
X"0177",
X"F7B3",
X"FAA1",
X"FE0C",
X"FD12",
X"FD8F",
X"FC18",
X"FB9B",
X"FC95",
X"F8AD",
X"FB9B",
X"F5BF",
X"F542",
X"EFE3",
X"ED72",
X"EBFB",
X"EA84",
X"EB01",
X"EB01",
X"EB7E",
X"EE6C",
X"EB01",
X"E90D",
X"E69C",
X"EBFB",
X"EFE3",
X"ECF5",
X"ECF5",
X"ED72",
X"EC78",
X"EF66",
X"F060",
X"ED72",
X"EDEF",
X"EF66",
X"EFE3",
X"EE6C",
X"F63C",
X"F34E",
X"F830",
X"FF06",
X"FB9B",
X"F8AD",
X"F736",
X"03E8",
X"007D",
X"0465",
X"0465",
X"02EE",
X"02EE",
X"0465",
X"FF83",
X"0177",
X"0177",
X"007D",
X"036B",
X"0753",
X"02EE",
X"05DC",
X"05DC",
X"0465",
X"007D",
X"FAA1",
X"03E8",
X"055F",
X"03E8",
X"0271",
X"036B",
X"0465",
X"09C4",
X"0659",
X"0947",
X"08CA",
X"055F",
X"04E2",
X"08CA",
X"03E8",
X"036B",
X"036B",
X"01F4",
X"0271",
X"03E8",
X"03E8",
X"FE0C",
X"FA24",
X"FB9B",
X"FD8F",
X"FE89",
X"F63C",
X"FAA1",
X"F5BF",
X"F63C",
X"F6B9",
X"F5BF",
X"FE89",
X"F542",
X"FD12",
X"036B",
X"FD12",
X"FF06",
X"0659",
X"0D2F",
X"0177",
X"07D0",
X"0753",
X"0BB8",
X"0FA0",
X"0FA0",
X"1117",
X"101D",
X"0DAC",
X"0EA6",
X"128E",
X"1388",
X"128E",
X"0D2F",
X"06D6",
X"0753",
X"06D6",
X"084D",
X"0BB8",
X"0ABE",
X"07D0",
X"06D6",
X"055F",
X"0271",
X"084D",
X"05DC",
X"0D2F",
X"0E29",
X"09C4",
X"0C35",
X"0DAC",
X"09C4",
X"0FA0",
X"0F23",
X"0F23",
X"0D2F",
X"109A",
X"15F9",
X"0DAC",
X"14FF",
X"101D",
X"0FA0",
X"0B3B",
X"06D6",
X"04E2",
X"055F",
X"0659",
X"00FA",
X"0947",
X"0F23",
X"0ABE",
X"0A41",
X"0C35",
X"0947",
X"0947",
X"07D0",
X"0659",
X"055F",
X"0271",
X"036B",
X"084D",
X"0C35",
X"0D2F",
X"0753",
X"09C4",
X"00FA",
X"FE0C",
X"FF83",
X"FB1E",
X"FB1E",
X"F8AD",
X"F5BF",
X"FAA1",
X"007D",
X"007D",
X"FE89",
X"FD12",
X"FD12",
X"FE0C",
X"0177",
X"FA24",
X"FA24",
X"F8AD",
X"F5BF",
X"F2D1",
X"F63C",
X"F5BF",
X"F3CB",
X"EFE3",
X"F2D1",
X"F7B3",
X"F736",
X"F254",
X"F060",
X"F34E",
X"F448",
X"F6B9",
X"FA24",
X"F830",
X"FB9B",
X"FB9B",
X"007D",
X"F736",
X"FB1E",
X"FF06",
X"F542",
X"F5BF",
X"F6B9",
X"F542",
X"F5BF",
X"EFE3",
X"EE6C",
X"F2D1",
X"EF66",
X"ECF5",
X"E813",
X"ECF5",
X"E90D",
X"ED72",
X"EB7E",
X"E796",
X"E890",
X"EA07",
X"E813",
X"E796",
X"EB7E",
X"ECF5",
X"ECF5",
X"E796",
X"EA07",
X"E719",
X"EC78",
X"EF66",
X"EB01",
X"EB7E",
X"ED72",
X"EA84",
X"E4A8",
X"E813",
X"E3AE",
X"E2B4",
X"E331",
X"DDD2",
X"D9EA",
X"DCD8",
X"E61F",
X"E813",
X"E90D",
X"E890",
X"ECF5",
X"ED72",
X"EDEF",
X"EA07",
X"EB7E",
X"F1D7",
X"E813",
X"E813",
X"E42B",
X"E796",
X"E525",
X"E719",
X"E69C",
X"E331",
X"EA07",
X"E90D",
X"F2D1",
X"F5BF",
X"FB9B",
X"FD12",
X"FA24",
X"FD8F",
X"06D6",
X"04E2",
X"0753",
X"084D",
X"0271",
X"00FA",
X"FF06",
X"0177",
X"0659",
X"0F23",
X"0BB8",
X"128E",
X"1117",
X"1194",
X"128E",
X"109A",
X"130B",
X"130B",
X"17ED",
X"15F9",
X"1964",
X"1D4C",
X"1CCF",
X"1F40",
X"280A",
X"2134",
X"249F",
X"2981",
X"20B7",
X"2616",
X"23A5",
X"23A5",
X"1F40",
X"21B1",
X"1EC3",
X"1B58",
X"2134",
X"17ED",
X"1211",
X"1676",
X"109A",
X"130B",
X"1194",
X"0F23",
X"0EA6",
X"0DAC",
X"0CB2",
X"0C35",
X"0947",
X"06D6",
X"03E8",
X"0177",
X"07D0",
X"0947",
X"00FA",
X"04E2",
X"0000",
X"055F",
X"06D6",
X"0C35",
X"0B3B",
X"0947",
X"0271",
X"0465",
X"02EE",
X"01F4",
X"0B3B",
X"007D",
X"05DC",
X"0BB8",
X"07D0",
X"09C4",
X"07D0",
X"07D0",
X"05DC",
X"06D6",
X"02EE",
X"03E8",
X"05DC",
X"FF06",
X"F8AD",
X"FD12",
X"FD12",
X"FC18",
X"FB1E",
X"F7B3",
X"FC18",
X"F9A7",
X"FD8F",
X"FD12",
X"FF83",
X"036B",
X"02EE",
X"084D",
X"0753",
X"05DC",
X"036B",
X"08CA",
X"0659",
X"055F",
X"06D6",
X"07D0",
X"04E2",
X"01F4",
X"04E2",
X"06D6",
X"0D2F",
X"0CB2",
X"1482",
X"0B3B",
X"09C4",
X"055F",
X"02EE",
X"09C4",
X"04E2",
X"01F4",
X"04E2",
X"07D0",
X"0BB8",
X"0ABE",
X"09C4",
X"0CB2",
X"0753",
X"05DC",
X"04E2",
X"0659",
X"0659",
X"036B",
X"0947",
X"0177",
X"FE89",
X"02EE",
X"036B",
X"FE0C",
X"FE89",
X"FE89",
X"007D",
X"0465",
X"FC95",
X"FB9B",
X"00FA",
X"FB9B",
X"FD8F",
X"F9A7",
X"FC18",
X"FD12",
X"0177",
X"03E8",
X"FE89",
X"FF83",
X"FC95",
X"00FA",
X"01F4",
X"00FA",
X"FE89",
X"F9A7",
X"FF06",
X"0000",
X"0000",
X"FC95",
X"FB1E",
X"00FA",
X"01F4",
X"0465",
X"02EE",
X"0753",
X"0ABE",
X"07D0",
X"0B3B",
X"00FA",
X"04E2",
X"FF83",
X"FB9B",
X"036B",
X"FA24",
X"FC95",
X"0177",
X"055F",
X"036B",
X"FF83",
X"00FA",
X"FE89",
X"0000",
X"04E2",
X"FE89",
X"FD8F",
X"00FA",
X"FA24",
X"FC18",
X"FF83",
X"0465",
X"0BB8",
X"05DC",
X"04E2",
X"FB9B",
X"FC18",
X"FAA1",
X"F5BF",
X"F830",
X"F736",
X"FAA1",
X"FC95",
X"F92A",
X"F7B3",
X"007D",
X"FE0C",
X"F542",
X"F8AD",
X"F254",
X"F3CB",
X"F6B9",
X"F5BF",
X"F5BF",
X"F6B9",
X"F1D7",
X"F4C5",
X"F254",
X"EF66",
X"EE6C",
X"F34E",
X"F4C5",
X"F3CB",
X"F448",
X"F0DD",
X"F3CB",
X"F34E",
X"EF66",
X"F1D7",
X"F0DD",
X"E98A",
X"E719",
X"F2D1",
X"EFE3",
X"EFE3",
X"F9A7",
X"F4C5",
X"F63C",
X"FA24",
X"F5BF",
X"F3CB",
X"F736",
X"F63C",
X"F1D7",
X"F542",
X"F254",
X"F254",
X"F736",
X"F3CB",
X"EFE3",
X"F15A",
X"F34E",
X"F6B9",
X"F0DD",
X"ED72",
X"F34E",
X"F060",
X"F6B9",
X"F63C",
X"FE0C",
X"06D6",
X"00FA",
X"02EE",
X"03E8",
X"F8AD",
X"FC18",
X"FF83",
X"FD8F",
X"02EE",
X"FF83",
X"FB9B",
X"FC18",
X"01F4",
X"0000",
X"FE0C",
X"0000",
X"F8AD",
X"FB9B",
X"FAA1",
X"FE0C",
X"00FA",
X"0177",
X"0177",
X"055F",
X"03E8",
X"02EE",
X"055F",
X"04E2",
X"07D0",
X"036B",
X"0BB8",
X"08CA",
X"0B3B",
X"101D",
X"0465",
X"0947",
X"0ABE",
X"0753",
X"0ABE",
X"0753",
X"084D",
X"0947",
X"09C4",
X"0DAC",
X"0DAC",
X"1117",
X"1405",
X"09C4",
X"0D2F",
X"0EA6",
X"06D6",
X"FC18",
X"0177",
X"084D",
X"03E8",
X"03E8",
X"02EE",
X"04E2",
X"05DC",
X"05DC",
X"09C4",
X"04E2",
X"0177",
X"FE89",
X"FE0C",
X"FD12",
X"F9A7",
X"F63C",
X"FC95",
X"FC95",
X"FAA1",
X"F830",
X"F9A7",
X"FF83",
X"FAA1",
X"FC95",
X"084D",
X"FF06",
X"0A41",
X"08CA",
X"FD8F",
X"04E2",
X"07D0",
X"FD8F",
X"FB1E",
X"F736",
X"F34E",
X"F34E",
X"ECF5",
X"F542",
X"F6B9",
X"F5BF",
X"007D",
X"FA24",
X"00FA",
X"09C4",
X"01F4",
X"02EE",
X"0A41",
X"08CA",
X"06D6",
X"101D",
X"0C35",
X"1117",
X"1117",
X"1117",
X"130B",
X"109A",
X"0A41",
X"055F",
X"0BB8",
X"036B",
X"0ABE",
X"0465",
X"FD12",
X"07D0",
X"0465",
X"0B3B",
X"00FA",
X"06D6",
X"007D",
X"FD8F",
X"0DAC",
X"02EE",
X"055F",
X"00FA",
X"F6B9",
X"FE89",
X"F4C5",
X"F830",
X"F1D7",
X"F060",
X"F4C5",
X"ED72",
X"F254",
X"EDEF",
X"F1D7",
X"EE6C",
X"F63C",
X"FC18",
X"EFE3",
X"F4C5",
X"F0DD",
X"F9A7",
X"F92A",
X"EFE3",
X"F63C",
X"F542",
X"F34E",
X"F060",
X"F254",
X"F34E",
X"FA24",
X"007D",
X"02EE",
X"06D6",
X"036B",
X"01F4",
X"03E8",
X"0753",
X"01F4",
X"055F",
X"0659",
X"07D0",
X"0947",
X"0ABE",
X"09C4",
X"07D0",
X"0D2F",
X"0E29",
X"0ABE",
X"0C35",
X"109A",
X"1676",
X"19E1",
X"1964",
X"1B58",
X"1770",
X"1770",
X"1482",
X"1482",
X"1C52",
X"19E1",
X"1EC3",
X"1ADB",
X"1117",
X"109A",
X"130B",
X"0DAC",
X"0271",
X"07D0",
X"09C4",
X"0465",
X"07D0",
X"08CA",
X"07D0",
X"0659",
X"FC95",
X"00FA",
X"FB9B",
X"FD8F",
X"FAA1",
X"F9A7",
X"F254",
X"F830",
X"FC95",
X"F736",
X"0271",
X"FC95",
X"FD8F",
X"FAA1",
X"F2D1",
X"F254",
X"F060",
X"EFE3",
X"F060",
X"F254",
X"EBFB",
X"EC78",
X"E3AE",
X"E043",
X"E42B",
X"DECC",
X"E2B4",
X"E13D",
X"DECC",
X"E813",
X"EFE3",
X"EFE3",
X"ECF5",
X"F1D7",
X"EF66",
X"EA07",
X"ED72",
X"EA07",
X"EB7E",
X"E98A",
X"ED72",
X"E813",
X"E0C0",
X"DFC6",
X"DECC",
X"E69C",
X"E331",
X"E69C",
X"EFE3",
X"E90D",
X"EB7E",
X"F0DD",
X"ECF5",
X"EFE3",
X"F254",
X"F2D1",
X"EEE9",
X"F34E",
X"F3CB",
X"F3CB",
X"F6B9",
X"F448",
X"F448",
X"EB01",
X"EBFB",
X"F3CB",
X"F254",
X"FB1E",
X"FD8F",
X"F9A7",
X"FB9B",
X"F92A",
X"FB1E",
X"007D",
X"04E2",
X"0465",
X"06D6",
X"0271",
X"00FA",
X"00FA",
X"007D",
X"03E8",
X"09C4",
X"0E29",
X"0947",
X"0EA6",
X"1405",
X"0C35",
X"07D0",
X"08CA",
X"0753",
X"0000",
X"FE89",
X"084D",
X"0FA0",
X"0FA0",
X"1194",
X"1770",
X"130B",
X"1770",
X"15F9",
X"14FF",
X"1B58",
X"1405",
X"1211",
X"1194",
X"101D",
X"0F23",
X"0FA0",
X"1405",
X"1482",
X"0EA6",
X"14FF",
X"1388",
X"1482",
X"15F9",
X"1770",
X"1F40",
X"18E7",
X"1770",
X"1676",
X"1482",
X"16F3",
X"19E1",
X"1964",
X"1676",
X"17ED",
X"1405",
X"186A",
X"1770",
X"1770",
X"1A5E",
X"1D4C",
X"1EC3",
X"1BD5",
X"16F3",
X"1676",
X"18E7",
X"18E7",
X"130B",
X"1211",
X"0EA6",
X"1388",
X"109A",
X"128E",
X"1676",
X"0F23",
X"1388",
X"1ADB",
X"1A5E",
X"1BD5",
X"203A",
X"186A",
X"2422",
X"18E7",
X"128E",
X"0E29",
X"0C35",
X"0FA0",
X"0E29",
X"157C",
X"186A",
X"2328",
X"2422",
X"2904",
X"2693",
X"280A",
X"278D",
X"1F40",
X"1A5E",
X"1388",
X"0753",
X"0947",
X"FD8F",
X"01F4",
X"0BB8",
X"007D",
X"0177",
X"06D6",
X"0C35",
X"03E8",
X"04E2",
X"0177",
X"055F",
X"0271",
X"0000",
X"FB9B",
X"FE0C",
X"036B",
X"0000",
X"0271",
X"FE0C",
X"FD12",
X"03E8",
X"036B",
X"FD12",
X"007D",
X"F92A",
X"0000",
X"F1D7",
X"EA84",
X"E2B4",
X"E4A8",
X"DFC6",
X"DFC6",
X"E331",
X"DBDE",
X"D585",
X"D21A",
X"D67F",
X"DA67",
X"DB61",
X"DF49",
X"DFC6",
X"DCD8",
X"DC5B",
X"D96D",
X"D508",
X"D297",
X"D026",
X"CF2C",
X"D585",
X"D391",
X"D314",
X"D0A3",
X"D120",
X"CDB5",
X"CFA9",
X"D026",
X"D19D",
X"D67F",
X"D391",
X"D48B",
X"D120",
X"CFA9",
X"D391",
X"D297",
X"D120",
X"CFA9",
X"CA4A",
X"CCBB",
X"D026",
X"D0A3",
X"D40E",
X"D508",
X"D873",
X"DECC",
X"D9EA",
X"DF49",
X"E043",
X"DC5B",
X"DECC",
X"DA67",
X"D602",
X"D779",
X"D67F",
X"DD55",
X"E331",
X"DECC",
X"DC5B",
X"DBDE",
X"E3AE",
X"E796",
X"EA07",
X"E90D",
X"E890",
X"EBFB",
X"EDEF",
X"F0DD",
X"F7B3",
X"FC18",
X"FAA1",
X"FE89",
X"FB9B",
X"FB1E",
X"FB1E",
X"F736",
X"F92A",
X"FD12",
X"FB9B",
X"FC95",
X"FF83",
X"FF83",
X"FC95",
X"00FA",
X"01F4",
X"07D0",
X"0D2F",
X"0E29",
X"0F23",
X"128E",
X"130B",
X"1405",
X"0E29",
X"0F23",
X"1194",
X"1388",
X"1117",
X"186A",
X"16F3",
X"186A",
X"2134",
X"22AB",
X"29FE",
X"2616",
X"2E63",
X"29FE",
X"30D4",
X"2F5D",
X"2616",
X"2C6F",
X"2981",
X"2E63",
X"3057",
X"2D69",
X"2616",
X"2422",
X"2616",
X"21B1",
X"2134",
X"20B7",
X"1CCF",
X"1DC9",
X"203A",
X"2422",
X"22AB",
X"23A5",
X"1D4C",
X"1F40",
X"1F40",
X"1770",
X"17ED",
X"18E7",
X"17ED",
X"14FF",
X"1964",
X"1B58",
X"1ADB",
X"1BD5",
X"203A",
X"1B58",
X"1482",
X"1405",
X"128E",
X"1117",
X"0D2F",
X"09C4",
X"0465",
X"0947",
X"16F3",
X"1194",
X"130B",
X"1211",
X"1194",
X"0C35",
X"0947",
X"04E2",
X"0947",
X"02EE",
X"FD12",
X"007D",
X"0000",
X"04E2",
X"0A41",
X"0A41",
X"084D",
X"0753",
X"007D",
X"0177",
X"06D6",
X"0000",
X"FC18",
X"01F4",
X"FF83",
X"FB9B",
X"007D",
X"FB9B",
X"F9A7",
X"FE89",
X"0465",
X"FF83",
X"084D",
X"0CB2",
X"0D2F",
X"101D",
X"0ABE",
X"0C35",
X"0DAC",
X"06D6",
X"0BB8",
X"09C4",
X"0753",
X"0ABE",
X"0EA6",
X"08CA",
X"0659",
X"0ABE",
X"055F",
X"0753",
X"09C4",
X"07D0",
X"055F",
X"055F",
X"00FA",
X"055F",
X"0947",
X"0ABE",
X"084D",
X"05DC",
X"FF83",
X"FF83",
X"06D6",
X"FF06",
X"0177",
X"F9A7",
X"ED72",
X"E98A",
X"EC78",
X"ECF5",
X"EA07",
X"EB01",
X"EA84",
X"EE6C",
X"F3CB",
X"F2D1",
X"F254",
X"F254",
X"EFE3",
X"ED72",
X"E69C",
X"E5A2",
X"E4A8",
X"E42B",
X"E69C",
X"E2B4",
X"DF49",
X"DAE4",
X"DE4F",
X"E043",
X"E043",
X"E3AE",
X"E13D",
X"DFC6",
X"E813",
X"EE6C",
X"ECF5",
X"F34E",
X"EEE9",
X"F736",
X"FAA1",
X"F542",
X"F63C",
X"F2D1",
X"F1D7",
X"F15A",
X"F3CB",
X"F3CB",
X"F7B3",
X"F6B9",
X"FB9B",
X"FB9B",
X"00FA",
X"0465",
X"007D",
X"007D",
X"FD12",
X"0271",
X"FF06",
X"F7B3",
X"F736",
X"FD12",
X"F9A7",
X"FAA1",
X"0271",
X"FAA1",
X"FF06",
X"0271",
X"0000",
X"01F4",
X"05DC",
X"0753",
X"0753",
X"05DC",
X"0B3B",
X"0947",
X"01F4",
X"03E8",
X"04E2",
X"03E8",
X"FD8F",
X"0177",
X"05DC",
X"FF06",
X"036B",
X"FF06",
X"04E2",
X"05DC",
X"03E8",
X"00FA",
X"03E8",
X"0947",
X"007D",
X"036B",
X"FE0C",
X"01F4",
X"08CA",
X"00FA",
X"01F4",
X"01F4",
X"00FA",
X"03E8",
X"01F4",
X"F8AD",
X"F8AD",
X"FD8F",
X"FB9B",
X"FC18",
X"01F4",
X"FE89",
X"05DC",
X"0EA6",
X"1194",
X"0DAC",
X"1388",
X"0F23",
X"055F",
X"036B",
X"0000",
X"FE89",
X"FD8F",
X"F3CB",
X"F254",
X"EE6C",
X"EBFB",
X"ECF5",
X"ED72",
X"F5BF",
X"FAA1",
X"F5BF",
X"FAA1",
X"F92A",
X"FC95",
X"FD8F",
X"FC18",
X"007D",
X"0000",
X"FB1E",
X"007D",
X"0465",
X"0659",
X"0947",
X"06D6",
X"08CA",
X"0D2F",
X"0A41",
X"0A41",
X"0EA6",
X"0C35",
X"0753",
X"04E2",
X"055F",
X"04E2",
X"0A41",
X"06D6",
X"0177",
X"05DC",
X"0465",
X"0CB2",
X"0B3B",
X"03E8",
X"08CA",
X"0B3B",
X"0F23",
X"0F23",
X"0FA0",
X"0EA6",
X"0B3B",
X"109A",
X"101D",
X"0FA0",
X"109A",
X"0EA6",
X"0C35",
X"0947",
X"0F23",
X"1211",
X"0CB2",
X"084D",
X"06D6",
X"0947",
X"08CA",
X"0BB8",
X"0B3B",
X"FB9B",
X"0271",
X"02EE",
X"02EE",
X"03E8",
X"FE0C",
X"0753",
X"0ABE",
X"0ABE",
X"0C35",
X"09C4",
X"0C35",
X"084D",
X"04E2",
X"FE89",
X"F830",
X"FB1E",
X"F6B9",
X"EEE9",
X"EE6C",
X"EB7E",
X"ECF5",
X"ECF5",
X"EEE9",
X"ED72",
X"EFE3",
X"EA07",
X"E5A2",
X"E719",
X"E1BA",
X"DDD2",
X"DCD8",
X"DDD2",
X"E890",
X"E890",
X"E69C",
X"E1BA",
X"E69C",
X"ED72",
X"EDEF",
X"ED72",
X"EBFB",
X"EA84",
X"EC78",
X"E796",
X"E5A2",
X"E813",
X"EA84",
X"EFE3",
X"F3CB",
X"F2D1",
X"F1D7",
X"F1D7",
X"F1D7",
X"F5BF",
X"F8AD",
X"F736",
X"F5BF",
X"F736",
X"FA24",
X"FC18",
X"FC18",
X"0271",
X"01F4",
X"FE0C",
X"0000",
X"FC95",
X"055F",
X"0465",
X"05DC",
X"05DC",
X"055F",
X"03E8",
X"0000",
X"FC95",
X"F34E",
X"F34E",
X"EFE3",
X"F060",
X"E890",
X"E2B4",
X"E331",
X"E90D",
X"E890",
X"E98A",
X"E69C",
X"EA07",
X"ECF5",
X"EE6C",
X"EBFB",
X"EB7E",
X"EBFB",
X"EB7E",
X"EFE3",
X"F15A",
X"F830",
X"FD8F",
X"FD8F",
X"FC95",
X"F542",
X"FD12",
X"007D",
X"FAA1",
X"FC18",
X"F6B9",
X"F5BF",
X"FD12",
X"F830",
X"F8AD",
X"0000",
X"FC18",
X"0271",
X"055F",
X"055F",
X"0ABE",
X"0D2F",
X"128E",
X"14FF",
X"1117",
X"128E",
X"14FF",
X"109A",
X"1194",
X"1211",
X"1405",
X"1482",
X"1ADB",
X"2134",
X"2134",
X"2134",
X"1CCF",
X"1CCF",
X"19E1",
X"15F9",
X"1211",
X"101D",
X"109A",
X"1117",
X"1405",
X"186A",
X"1ADB",
X"1405",
X"1482",
X"157C",
X"18E7",
X"1EC3",
X"1E46",
X"21B1",
X"249F",
X"23A5",
X"249F",
X"249F",
X"249F",
X"2599",
X"278D",
X"2599",
X"2616",
X"2710",
X"2134",
X"2422",
X"1BD5",
X"1F40",
X"2328",
X"20B7",
X"2710",
X"1FBD",
X"21B1",
X"1D4C",
X"222E",
X"1CCF",
X"1B58",
X"1CCF",
X"1DC9",
X"15F9",
X"1388",
X"109A",
X"1117",
X"0CB2",
X"0EA6",
X"130B",
X"0947",
X"084D",
X"036B",
X"0177",
X"084D",
X"0659",
X"02EE",
X"05DC",
X"FD8F",
X"FE0C",
X"FF83",
X"F6B9",
X"F4C5",
X"F736",
X"F830",
X"F542",
X"F4C5",
X"FB1E",
X"FF06",
X"FD12",
X"FD8F",
X"036B",
X"0659",
X"0659",
X"0000",
X"FE0C",
X"02EE",
X"0659",
X"03E8",
X"03E8",
X"02EE",
X"05DC",
X"0659",
X"036B",
X"FD12",
X"007D",
X"FE89",
X"F830",
X"FB9B",
X"F3CB",
X"0271",
X"F9A7",
X"FA24",
X"0271",
X"0465",
X"036B",
X"0753",
X"08CA",
X"055F",
X"04E2",
X"0753",
X"07D0",
X"055F",
X"0BB8",
X"0177",
X"01F4",
X"06D6",
X"055F",
X"FC18",
X"F7B3",
X"FAA1",
X"FA24",
X"F3CB",
X"F3CB",
X"EC78",
X"E719",
X"EA84",
X"DFC6",
X"E4A8",
X"E42B",
X"E42B",
X"E237",
X"DFC6",
X"E043",
X"E4A8",
X"E0C0",
X"E237",
X"E2B4",
X"D9EA",
X"DDD2",
X"D508",
X"D602",
X"DFC6",
X"D21A",
X"D6FC",
X"D9EA",
X"D585",
X"D8F0",
X"D7F6",
X"DA67",
X"DE4F",
X"E42B",
X"EA07",
X"E890",
X"DECC",
X"E525",
X"E525",
X"E525",
X"E719",
X"E2B4",
X"E525",
X"DFC6",
X"DE4F",
X"DECC",
X"E69C",
X"D9EA",
X"DA67",
X"DECC",
X"DE4F",
X"E043",
X"E5A2",
X"E61F",
X"E525",
X"E796",
X"E331",
X"EB7E",
X"E90D",
X"E2B4",
X"E237",
X"E796",
X"EB01",
X"EEE9",
X"F7B3",
X"F736",
X"F542",
X"FB1E",
X"FE0C",
X"FF06",
X"04E2",
X"084D",
X"00FA",
X"0947",
X"FF06",
X"0BB8",
X"0947",
X"04E2",
X"0DAC",
X"055F",
X"0753",
X"0271",
X"007D",
X"FF83",
X"FE89",
X"FD8F",
X"FF83",
X"FE0C",
X"FB9B",
X"FD12",
X"FD12",
X"FD12",
X"FC95",
X"F5BF",
X"F2D1",
X"F736",
X"F254",
X"EB01",
X"E90D",
X"E90D",
X"EB7E",
X"E796",
X"EA07",
X"EDEF",
X"EB01",
X"E98A",
X"EFE3",
X"F3CB",
X"EEE9",
X"F448",
X"F060",
X"F34E",
X"F736",
X"F060",
X"F34E",
X"F7B3",
X"F8AD",
X"FE0C",
X"00FA",
X"03E8",
X"FF06",
X"06D6",
X"01F4",
X"0271",
X"04E2",
X"0659",
X"08CA",
X"0ABE",
X"0ABE",
X"0659",
X"0465",
X"0BB8",
X"08CA",
X"05DC",
X"109A",
X"0EA6",
X"0DAC",
X"0B3B",
X"1211",
X"1770",
X"0E29",
X"1194",
X"203A",
X"1B58",
X"157C",
X"1DC9",
X"2422",
X"23A5",
X"1D4C",
X"1FBD",
X"280A",
X"2DE6",
X"2981",
X"2887",
X"2D69",
X"33C2",
X"34BC",
X"33C2",
X"3151",
X"3057",
X"31CE",
X"3345",
X"343F",
X"33C2",
X"3057",
X"2EE0",
X"2EE0",
X"3539",
X"33C2",
X"2FDA",
X"343F",
X"2EE0",
X"29FE",
X"2BF2",
X"2CEC",
X"2BF2",
X"2A7B",
X"3057",
X"2E63",
X"2A7B",
X"2BF2",
X"23A5",
X"2422",
X"2693",
X"22AB",
X"20B7",
X"1DC9",
X"21B1",
X"20B7",
X"1BD5",
X"1676",
X"157C",
X"186A",
X"1117",
X"101D",
X"0CB2",
X"09C4",
X"09C4",
X"08CA",
X"0947",
X"05DC",
X"FF83",
X"FF06",
X"03E8",
X"084D",
X"00FA",
X"055F",
X"08CA",
X"FF83",
X"0177",
X"0ABE",
X"084D",
X"055F",
X"08CA",
X"09C4",
X"07D0",
X"03E8",
X"FE89",
X"03E8",
X"0DAC",
X"0000",
X"FD8F",
X"02EE",
X"FE0C",
X"F9A7",
X"FB9B",
X"F8AD",
X"EF66",
X"F2D1",
X"F542",
X"ED72",
X"E331",
X"DFC6",
X"E4A8",
X"E61F",
X"E525",
X"DE4F",
X"DB61",
X"D779",
X"DA67",
X"DD55",
X"DCD8",
X"D96D",
X"D9EA",
X"DCD8",
X"D602",
X"D602",
X"D602",
X"D585",
X"D67F",
X"D9EA",
X"DECC",
X"DDD2",
X"D508",
X"DDD2",
X"DAE4",
X"D48B",
X"D391",
X"D602",
X"D585",
X"D026",
X"D026",
X"D391",
X"D0A3",
X"D67F",
X"D391",
X"CE32",
X"CFA9",
X"D6FC",
X"D0A3",
X"DD55",
X"DAE4",
X"D602",
X"D21A",
X"DC5B",
X"DA67",
X"DE4F",
X"E2B4",
X"E1BA",
X"EA84",
X"E237",
X"E719",
X"EB01",
X"EA84",
X"F4C5",
X"F060",
X"F2D1",
X"F8AD",
X"EEE9",
X"F4C5",
X"F3CB",
X"F736",
X"EBFB",
X"F0DD",
X"F060",
X"F1D7",
X"F542",
X"EFE3",
X"F448",
X"F254",
X"F7B3",
X"F4C5",
X"F92A",
X"02EE",
X"FB9B",
X"FAA1",
X"FB9B",
X"036B",
X"FB1E",
X"FF83",
X"FAA1",
X"FC18",
X"007D",
X"FB1E",
X"0271",
X"FD12",
X"FAA1",
X"036B",
X"01F4",
X"02EE",
X"0947",
X"0B3B",
X"0271",
X"055F",
X"0271",
X"07D0",
X"0CB2",
X"0DAC",
X"0F23",
X"0DAC",
X"0F23",
X"0D2F",
X"0CB2",
X"0B3B",
X"0947",
X"109A",
X"1388",
X"1211",
X"0F23",
X"0FA0",
X"0A41",
X"109A",
X"1482",
X"0C35",
X"0B3B",
X"0B3B",
X"0CB2",
X"05DC",
X"1194",
X"1211",
X"1194",
X"0E29",
X"1211",
X"186A",
X"186A",
X"1EC3",
X"1CCF",
X"2422",
X"1EC3",
X"1F40",
X"2422",
X"278D",
X"2599",
X"2616",
X"2F5D",
X"2B75",
X"2981",
X"2D69",
X"2981",
X"278D",
X"29FE",
X"2599",
X"2599",
X"2134",
X"1D4C",
X"1C52",
X"1676",
X"1964",
X"17ED",
X"130B",
X"0C35",
X"0BB8",
X"0F23",
X"0C35",
X"0EA6",
X"08CA",
X"0465",
X"0271",
X"00FA",
X"036B",
X"007D",
X"01F4",
X"FB1E",
X"F254",
X"F1D7",
X"F34E",
X"F830",
X"F736",
X"EC78",
X"EDEF",
X"F830",
X"F3CB",
X"F34E",
X"F7B3",
X"F736",
X"F34E",
X"F4C5",
X"F254",
X"F254",
X"EE6C",
X"EB7E",
X"F2D1",
X"EB01",
X"EE6C",
X"EF66",
X"EDEF",
X"F1D7",
X"F34E",
X"F1D7",
X"F9A7",
X"F5BF",
X"F6B9",
X"F1D7",
X"F4C5",
X"FF06",
X"F5BF",
X"F542",
X"00FA",
X"00FA",
X"0177",
X"0000",
X"00FA",
X"FD8F",
X"FAA1",
X"00FA",
X"007D",
X"036B",
X"0D2F",
X"0DAC",
X"0A41",
X"0B3B",
X"0F23",
X"0659",
X"09C4",
X"0ABE",
X"0A41",
X"0ABE",
X"0DAC",
X"0FA0",
X"1117",
X"0CB2",
X"1388",
X"130B",
X"1A5E",
X"1B58",
X"1405",
X"1B58",
X"16F3",
X"15F9",
X"14FF",
X"1482",
X"17ED",
X"16F3",
X"157C",
X"157C",
X"18E7",
X"1ADB",
X"128E",
X"109A",
X"186A",
X"1B58",
X"15F9",
X"15F9",
X"1405",
X"101D",
X"0FA0",
X"0EA6",
X"0BB8",
X"0F23",
X"09C4",
X"0753",
X"0B3B",
X"08CA",
X"0465",
X"084D",
X"00FA",
X"007D",
X"01F4",
X"FF06",
X"FD12",
X"F7B3",
X"F448",
X"F060",
X"ED72",
X"EC78",
X"EB7E",
X"E331",
X"E331",
X"E813",
X"E13D",
X"E3AE",
X"E61F",
X"E1BA",
X"E1BA",
X"E3AE",
X"E42B",
X"DF49",
X"DECC",
X"E0C0",
X"E237",
X"E043",
X"E525",
X"E813",
X"E719",
X"E61F",
X"E90D",
X"EA07",
X"EB01",
X"E90D",
X"E525",
X"E61F",
X"EBFB",
X"EC78",
X"EDEF",
X"F0DD",
X"F3CB",
X"FAA1",
X"F92A",
X"F7B3",
X"FC18",
X"FD12",
X"02EE",
X"00FA",
X"02EE",
X"0465",
X"FE89",
X"FC95",
X"F736",
X"F448",
X"F542",
X"F3CB",
X"F1D7",
X"EF66",
X"ED72",
X"EEE9",
X"F2D1",
X"F1D7",
X"EE6C",
X"F2D1",
X"F060",
X"EB01",
X"F060",
X"EE6C",
X"EF66",
X"EF66",
X"ECF5",
X"EDEF",
X"EA07",
X"ED72",
X"ED72",
X"EB7E",
X"EA07",
X"E890",
X"E5A2",
X"E525",
X"E2B4",
X"E3AE",
X"E61F",
X"EB7E",
X"E813",
X"E61F",
X"EF66",
X"EE6C",
X"EEE9",
X"F448",
X"F63C",
X"EE6C",
X"EDEF",
X"F0DD",
X"EE6C",
X"F3CB",
X"F34E",
X"F448",
X"F3CB",
X"F92A",
X"FA24",
X"FC18",
X"FE0C",
X"F7B3",
X"FC18",
X"F92A",
X"FC95",
X"FD8F",
X"0271",
X"04E2",
X"0465",
X"0B3B",
X"04E2",
X"0659",
X"1194",
X"0EA6",
X"0E29",
X"101D",
X"130B",
X"157C",
X"1676",
X"186A",
X"186A",
X"1770",
X"1770",
X"1ADB",
X"1B58",
X"1676",
X"1405",
X"15F9",
X"157C",
X"1405",
X"1770",
X"157C",
X"1770",
X"15F9",
X"18E7",
X"19E1",
X"1DC9",
X"2134",
X"1E46",
X"2134",
X"1C52",
X"1CCF",
X"1EC3",
X"1F40",
X"1EC3",
X"1F40",
X"1FBD",
X"1A5E",
X"1DC9",
X"1DC9",
X"1CCF",
X"1ADB",
X"1C52",
X"1CCF",
X"1BD5",
X"1A5E",
X"1A5E",
X"1ADB",
X"19E1",
X"17ED",
X"186A",
X"1676",
X"1388",
X"1676",
X"1211",
X"128E",
X"128E",
X"1211",
X"0ABE",
X"055F",
X"08CA",
X"0C35",
X"0753",
X"02EE",
X"02EE",
X"0271",
X"02EE",
X"FD8F",
X"FD8F",
X"FE89",
X"F9A7",
X"FAA1",
X"FD8F",
X"FB9B",
X"F63C",
X"F736",
X"FA24",
X"F9A7",
X"F830",
X"FB1E",
X"FD8F",
X"F8AD",
X"007D",
X"0000",
X"0000",
X"0000",
X"0271",
X"055F",
X"0271",
X"03E8",
X"0753",
X"09C4",
X"0BB8",
X"08CA",
X"084D",
X"0A41",
X"0ABE",
X"0E29",
X"1117",
X"128E",
X"109A",
X"157C",
X"17ED",
X"130B",
X"1482",
X"1482",
X"1211",
X"0C35",
X"1676",
X"157C",
X"0C35",
X"14FF",
X"1405",
X"0E29",
X"0A41",
X"084D",
X"0A41",
X"05DC",
X"03E8",
X"0465",
X"0000",
X"036B",
X"FE89",
X"FF83",
X"0000",
X"0000",
X"FE89",
X"F7B3",
X"F9A7",
X"F8AD",
X"F6B9",
X"F2D1",
X"F0DD",
X"EE6C",
X"EE6C",
X"EDEF",
X"E813",
X"E813",
X"E90D",
X"EDEF",
X"E525",
X"E890",
X"E61F",
X"E2B4",
X"E42B",
X"E13D",
X"E1BA",
X"E813",
X"E890",
X"E69C",
X"EC78",
X"EA84",
X"EBFB",
X"ECF5",
X"E90D",
X"EB7E",
X"ED72",
X"EDEF",
X"EA84",
X"EC78",
X"ED72",
X"EB7E",
X"F0DD",
X"F15A",
X"F0DD",
X"F1D7",
X"F2D1",
X"F060",
X"F254",
X"F1D7",
X"F254",
X"F254",
X"EEE9",
X"EC78",
X"ECF5",
X"E90D",
X"EA84",
X"F254",
X"ED72",
X"E98A",
X"EFE3",
X"EEE9",
X"E90D",
X"EEE9",
X"F15A",
X"EA07",
X"F254",
X"EFE3",
X"F3CB",
X"F34E",
X"F736",
X"F7B3",
X"F2D1",
X"F830",
X"EFE3",
X"F448",
X"F63C",
X"F448",
X"FF06",
X"FF06",
X"F7B3",
X"FB9B",
X"FF06",
X"00FA",
X"007D",
X"055F",
X"05DC",
X"036B",
X"03E8",
X"00FA",
X"084D",
X"07D0",
X"0753",
X"09C4",
X"0A41",
X"0CB2",
X"0B3B",
X"04E2",
X"0465",
X"0947",
X"08CA",
X"08CA",
X"084D",
X"05DC",
X"06D6",
X"00FA",
X"0659",
X"04E2",
X"FF06",
X"FE0C",
X"FF06",
X"FAA1",
X"0177",
X"FAA1",
X"FD8F",
X"0000",
X"F9A7",
X"F9A7",
X"F5BF",
X"F8AD",
X"FB1E",
X"FB1E",
X"F34E",
X"F5BF",
X"FC95",
X"F6B9",
X"F448",
X"F5BF",
X"F830",
X"FB1E",
X"FAA1",
X"FC95",
X"FE89",
X"FB1E",
X"FF83",
X"05DC",
X"0000",
X"FD8F",
X"03E8",
X"0947",
X"04E2",
X"05DC",
X"0F23",
X"1211",
X"128E",
X"0ABE",
X"0E29",
X"1194",
X"14FF",
X"101D",
X"1405",
X"16F3",
X"109A",
X"1194",
X"16F3",
X"14FF",
X"128E",
X"130B",
X"0DAC",
X"1117",
X"15F9",
X"1770",
X"109A",
X"0DAC",
X"1211",
X"130B",
X"0DAC",
X"0FA0",
X"1194",
X"101D",
X"101D",
X"0DAC",
X"0DAC",
X"0B3B",
X"08CA",
X"084D",
X"0C35",
X"0CB2",
X"08CA",
X"0659",
X"06D6",
X"0659",
X"0ABE",
X"0B3B",
X"01F4",
X"07D0",
X"09C4",
X"08CA",
X"04E2",
X"0465",
X"07D0",
X"FF06",
X"FF06",
X"FAA1",
X"F830",
X"FD12",
X"FC18",
X"F92A",
X"FC95",
X"F9A7",
X"F8AD",
X"FAA1",
X"F9A7",
X"F92A",
X"F736",
X"F4C5",
X"F2D1",
X"F830",
X"F8AD",
X"F34E",
X"F6B9",
X"F34E",
X"F15A",
X"EEE9",
X"EF66",
X"EFE3",
X"EDEF",
X"EC78",
X"ECF5",
X"EDEF",
X"E98A",
X"E813",
X"EB7E",
X"EB7E",
X"E90D",
X"EA84",
X"EA07",
X"EA07",
X"E890",
X"E61F",
X"E525",
X"E331",
X"E813",
X"E719",
X"E69C",
X"E719",
X"E4A8",
X"EA84",
X"EC78",
X"EB01",
X"EFE3",
X"F2D1",
X"F254",
X"F448",
X"F736",
X"F92A",
X"FAA1",
X"FD8F",
X"FD8F",
X"0177",
X"0271",
X"05DC",
X"05DC",
X"08CA",
X"0947",
X"0CB2",
X"1117",
X"1676",
X"1964",
X"1A5E",
X"1A5E",
X"1A5E",
X"1C52",
X"1F40",
X"203A",
X"1FBD",
X"21B1",
X"2599",
X"2422",
X"2693",
X"2710",
X"249F",
X"2693",
X"249F",
X"2693",
X"251C",
X"222E",
X"249F",
X"2422",
X"249F",
X"20B7",
X"2693",
X"2134",
X"1DC9",
X"20B7",
X"1CCF",
X"1D4C",
X"20B7",
X"1DC9",
X"1CCF",
X"1ADB",
X"1BD5",
X"186A",
X"1405",
X"109A",
X"0E29",
X"0CB2",
X"09C4",
X"08CA",
X"0C35",
X"02EE",
X"06D6",
X"0753",
X"03E8",
X"03E8",
X"03E8",
X"007D",
X"FF83",
X"FE89",
X"F830",
X"0271",
X"F92A",
X"F7B3",
X"F6B9",
X"F4C5",
X"F6B9",
X"F542",
X"F736",
X"EE6C",
X"EF66",
X"F63C",
X"F2D1",
X"F4C5",
X"F3CB",
X"FAA1",
X"FA24",
X"FA24",
X"F6B9",
X"F92A",
X"FB9B",
X"F6B9",
X"F4C5",
X"F448",
X"F7B3",
X"F736",
X"F542",
X"F3CB",
X"F6B9",
X"F830",
X"F63C",
X"F4C5",
X"F448",
X"F5BF",
X"F63C",
X"F3CB",
X"F92A",
X"FAA1",
X"F7B3",
X"F9A7",
X"FC18",
X"FE89",
X"FC95",
X"F63C",
X"FAA1",
X"FD12",
X"FC18",
X"FB9B",
X"F6B9",
X"F830",
X"F4C5",
X"F1D7",
X"F15A",
X"EFE3",
X"EEE9",
X"EB01",
X"EB01",
X"F0DD",
X"ED72",
X"EFE3",
X"EF66",
X"EF66",
X"F34E",
X"E98A",
X"EDEF",
X"ED72",
X"ECF5",
X"EF66",
X"EDEF",
X"F34E",
X"F1D7",
X"ECF5",
X"EFE3",
X"F34E",
X"F15A",
X"F2D1",
X"F63C",
X"F060",
X"F34E",
X"F4C5",
X"F1D7",
X"EF66",
X"ECF5",
X"ECF5",
X"EEE9",
X"EB01",
X"E98A",
X"EDEF",
X"ED72",
X"EB01",
X"E813",
X"EA84",
X"ED72",
X"EB7E",
X"E813",
X"E90D",
X"EA07",
X"E69C",
X"E69C",
X"E3AE",
X"DF49",
X"E331",
X"E237",
X"E0C0",
X"DF49",
X"E2B4",
X"E890",
X"E525",
X"E719",
X"E890",
X"E796",
X"E98A",
X"E90D",
X"EBFB",
X"EB7E",
X"EBFB",
X"EDEF",
X"EFE3",
X"EF66",
X"F63C",
X"F6B9",
X"F9A7",
X"FC95",
X"FB1E",
X"FF83",
X"FF06",
X"FD12",
X"FF83",
X"00FA",
X"02EE",
X"036B",
X"0A41",
X"0B3B",
X"0EA6",
X"101D",
X"0E29",
X"1211",
X"1194",
X"128E",
X"0CB2",
X"0DAC",
X"0D2F",
X"0659",
X"036B",
X"05DC",
X"0177",
X"055F",
X"0A41",
X"0947",
X"09C4",
X"0C35",
X"0EA6",
X"101D",
X"18E7",
X"19E1",
X"186A",
X"1964",
X"1770",
X"1C52",
X"1ADB",
X"1DC9",
X"18E7",
X"1194",
X"1482",
X"1405",
X"16F3",
X"109A",
X"14FF",
X"1E46",
X"1CCF",
X"1DC9",
X"2422",
X"1DC9",
X"17ED",
X"1E46",
X"186A",
X"128E",
X"1676",
X"109A",
X"1482",
X"19E1",
X"128E",
X"14FF",
X"16F3",
X"1964",
X"1B58",
X"1CCF",
X"1E46",
X"1CCF",
X"1BD5",
X"1BD5",
X"15F9",
X"1482",
X"186A",
X"1194",
X"1676",
X"130B",
X"0FA0",
X"0E29",
X"0EA6",
X"130B",
X"130B",
X"101D",
X"1676",
X"1ADB",
X"1964",
X"1964",
X"1482",
X"109A",
X"0DAC",
X"0DAC",
X"0DAC",
X"0DAC",
X"0D2F",
X"084D",
X"0A41",
X"0CB2",
X"0C35",
X"0F23",
X"0EA6",
X"0CB2",
X"0A41",
X"0FA0",
X"0753",
X"01F4",
X"0753",
X"03E8",
X"05DC",
X"06D6",
X"055F",
X"0271",
X"04E2",
X"0271",
X"FE89",
X"0177",
X"FE89",
X"00FA",
X"F9A7",
X"FAA1",
X"0000",
X"FE89",
X"0177",
X"FD8F",
X"036B",
X"007D",
X"FF83",
X"FE0C",
X"FB9B",
X"FC18",
X"0000",
X"FA24",
X"F6B9",
X"FD12",
X"FAA1",
X"F830",
X"F34E",
X"F0DD",
X"F3CB",
X"F15A",
X"F2D1",
X"F15A",
X"F448",
X"F4C5",
X"F34E",
X"F830",
X"F7B3",
X"F1D7",
X"EEE9",
X"F0DD",
X"EB01",
X"EA84",
X"F060",
X"F15A",
X"F34E",
X"F1D7",
X"F63C",
X"F830",
X"F2D1",
X"F542",
X"FB1E",
X"F736",
X"F34E",
X"F15A",
X"F830",
X"FAA1",
X"F2D1",
X"F448",
X"F3CB",
X"F542",
X"F448",
X"F0DD",
X"EEE9",
X"F0DD",
X"F060",
X"F34E",
X"F15A",
X"F0DD",
X"F1D7",
X"ED72",
X"EE6C",
X"ECF5",
X"EB7E",
X"E890",
X"E796",
X"EA07",
X"E98A",
X"EA07",
X"E69C",
X"E813",
X"EB01",
X"EA84",
X"ED72",
X"F3CB",
X"F2D1",
X"F1D7",
X"F63C",
X"F4C5",
X"F7B3",
X"F6B9",
X"F92A",
X"FC95",
X"FA24",
X"F92A",
X"FA24",
X"F63C",
X"F4C5",
X"F34E",
X"F542",
X"F34E",
X"F1D7",
X"EFE3",
X"EFE3",
X"EF66",
X"F15A",
X"F0DD",
X"ED72",
X"EC78",
X"EFE3",
X"F060",
X"E813",
X"E98A",
X"E98A",
X"E719",
X"ED72",
X"EFE3",
X"F0DD",
X"F92A",
X"F63C",
X"FD8F",
X"007D",
X"FD8F",
X"055F",
X"0947",
X"04E2",
X"0659",
X"09C4",
X"0947",
X"0EA6",
X"1117",
X"0CB2",
X"0EA6",
X"0DAC",
X"0E29",
X"0F23",
X"08CA",
X"0C35",
X"08CA",
X"0465",
X"0B3B",
X"09C4",
X"055F",
X"0947",
X"08CA",
X"06D6",
X"055F",
X"0000",
X"0271",
X"FF83",
X"FC18",
X"01F4",
X"FE89",
X"FF06",
X"02EE",
X"FD8F",
X"007D",
X"FF06",
X"FA24",
X"01F4",
X"F830",
X"FA24",
X"FC18",
X"FB9B",
X"F9A7",
X"FF06",
X"FF06",
X"007D",
X"0753",
X"055F",
X"05DC",
X"055F",
X"0A41",
X"0DAC",
X"1194",
X"1194",
X"0E29",
X"1405",
X"157C",
X"157C",
X"15F9",
X"157C",
X"1FBD",
X"1A5E",
X"16F3",
X"186A",
X"15F9",
X"1211",
X"186A",
X"15F9",
X"0F23",
X"1388",
X"0CB2",
X"0D2F",
X"0CB2",
X"06D6",
X"05DC",
X"0659",
X"03E8",
X"036B",
X"01F4",
X"0177",
X"FC18",
X"FC95",
X"F254",
X"F1D7",
X"FA24",
X"F6B9",
X"FA24",
X"F5BF",
X"EFE3",
X"F4C5",
X"FC95",
X"F4C5",
X"F4C5",
X"FD12",
X"F542",
X"F9A7",
X"FF83",
X"F736",
X"F6B9",
X"FD12",
X"FB9B",
X"F448",
X"F3CB",
X"F92A",
X"FC95",
X"F542",
X"F63C",
X"007D",
X"01F4",
X"0177",
X"036B",
X"01F4",
X"0271",
X"0753",
X"05DC",
X"0ABE",
X"0ABE",
X"0753",
X"055F",
X"00FA",
X"036B",
X"0659",
X"0753",
X"0659",
X"0DAC",
X"0EA6",
X"0B3B",
X"084D",
X"084D",
X"07D0",
X"0ABE",
X"0ABE",
X"05DC",
X"09C4",
X"09C4",
X"055F",
X"04E2",
X"084D",
X"07D0",
X"0465",
X"0177",
X"06D6",
X"0271",
X"01F4",
X"055F",
X"05DC",
X"0659",
X"0659",
X"0753",
X"07D0",
X"0271",
X"036B",
X"0465",
X"FC18",
X"FF06",
X"0000",
X"0000",
X"FE0C",
X"F8AD",
X"FB9B",
X"FD12",
X"FC18",
X"FB9B",
X"FB1E",
X"FD12",
X"007D",
X"02EE",
X"036B",
X"007D",
X"007D",
X"0947",
X"09C4",
X"0465",
X"0947",
X"08CA",
X"08CA",
X"084D",
X"084D",
X"0659",
X"FF06",
X"036B",
X"0465",
X"007D",
X"0000",
X"08CA",
X"0BB8",
X"0947",
X"08CA",
X"084D",
X"0659",
X"055F",
X"05DC",
X"0271",
X"08CA",
X"0A41",
X"FF06",
X"07D0",
X"0177",
X"007D",
X"FE89",
X"FC95",
X"0271",
X"03E8",
X"02EE",
X"FF83",
X"03E8",
X"0465",
X"02EE",
X"007D",
X"04E2",
X"0947",
X"05DC",
X"0753",
X"04E2",
X"03E8",
X"036B",
X"FF83",
X"01F4",
X"00FA",
X"F7B3",
X"FC95",
X"0000",
X"0000",
X"FF06",
X"00FA",
X"FF83",
X"FF06",
X"007D",
X"F830",
X"F8AD",
X"FD8F",
X"FC95",
X"F63C",
X"F9A7",
X"F63C",
X"F15A",
X"F34E",
X"EE6C",
X"EE6C",
X"F060",
X"F15A",
X"EFE3",
X"F0DD",
X"F1D7",
X"F254",
X"ECF5",
X"F0DD",
X"FE0C",
X"F0DD",
X"EFE3",
X"F34E",
X"F6B9",
X"F3CB",
X"F34E",
X"F4C5",
X"F3CB",
X"F736",
X"FE89",
X"0177",
X"FA24",
X"FA24",
X"F542",
X"F8AD",
X"FA24",
X"F92A",
X"FC95",
X"FC95",
X"FA24",
X"FAA1",
X"FAA1",
X"FE89",
X"00FA",
X"FC95",
X"007D",
X"FF83",
X"FE89",
X"FD12",
X"007D",
X"0271",
X"0271",
X"05DC",
X"0659",
X"0000",
X"FB1E",
X"02EE",
X"01F4",
X"FD8F",
X"036B",
X"02EE",
X"FF06",
X"0271",
X"036B",
X"0465",
X"0000",
X"FD12",
X"01F4",
X"FB9B",
X"FC95",
X"0271",
X"F9A7",
X"F5BF",
X"F3CB",
X"F7B3",
X"F1D7",
X"F448",
X"F3CB",
X"EB7E",
X"EE6C",
X"F254",
X"EEE9",
X"ECF5",
X"EB7E",
X"EEE9",
X"F2D1",
X"F0DD",
X"F1D7",
X"F0DD",
X"F060",
X"F060",
X"F060",
X"F1D7",
X"F060",
X"F1D7",
X"F0DD",
X"F34E",
X"F0DD",
X"EFE3",
X"F448",
X"F3CB",
X"F542",
X"F060",
X"F060",
X"EFE3",
X"EE6C",
X"EDEF",
X"EF66",
X"ECF5",
X"EA07",
X"EC78",
X"EB7E",
X"EE6C",
X"ECF5",
X"EBFB",
X"ECF5",
X"F1D7",
X"F2D1",
X"F5BF",
X"F63C",
X"F92A",
X"F9A7",
X"F736",
X"FB9B",
X"FA24",
X"F8AD",
X"FE89",
X"0000",
X"FE89",
X"0000",
X"02EE",
X"05DC",
X"0753",
X"0ABE",
X"0C35",
X"0B3B",
X"07D0",
X"0A41",
X"0B3B",
X"0B3B",
X"0A41",
X"07D0",
X"0A41",
X"0947",
X"09C4",
X"084D",
X"055F",
X"055F",
X"055F",
X"02EE",
X"04E2",
X"09C4",
X"07D0",
X"06D6",
X"05DC",
X"05DC",
X"07D0",
X"0ABE",
X"0D2F",
X"0F23",
X"0EA6",
X"0B3B",
X"0DAC",
X"0E29",
X"0A41",
X"0B3B",
X"0E29",
X"0DAC",
X"0FA0",
X"1194",
X"1482",
X"157C",
X"186A",
X"1D4C",
X"1DC9",
X"1FBD",
X"1CCF",
X"15F9",
X"17ED",
X"17ED",
X"1ADB",
X"1DC9",
X"1DC9",
X"1ADB",
X"1A5E",
X"1CCF",
X"1A5E",
X"186A",
X"1C52",
X"1DC9",
X"1B58",
X"1964",
X"1A5E",
X"18E7",
X"1A5E",
X"1964",
X"19E1",
X"19E1",
X"186A",
X"16F3",
X"1770",
X"1ADB",
X"1DC9",
X"2422",
X"222E",
X"1F40",
X"1F40",
X"21B1",
X"203A",
X"2134",
X"2134",
X"1DC9",
X"19E1",
X"15F9",
X"1676",
X"17ED",
X"128E",
X"1770",
X"1E46",
X"1C52",
X"186A",
X"1964",
X"14FF",
X"1117",
X"0FA0",
X"1482",
X"130B",
X"0FA0",
X"0EA6",
X"101D",
X"0D2F",
X"0CB2",
X"0DAC",
X"0E29",
X"0B3B",
X"0659",
X"06D6",
X"055F",
X"01F4",
X"FF06",
X"FAA1",
X"F63C",
X"F542",
X"F34E",
X"F254",
X"F448",
X"F5BF",
X"FAA1",
X"FF83",
X"FC18",
X"FAA1",
X"FD8F",
X"FC18",
X"F92A",
X"F34E",
X"ECF5",
X"EB01",
X"E719",
X"E237",
X"E3AE",
X"E42B",
X"E237",
X"E1BA",
X"DD55",
X"DF49",
X"E0C0",
X"E0C0",
X"E331",
X"E3AE",
X"EA07",
X"EB01",
X"E813",
X"E5A2",
X"E5A2",
X"E13D",
X"DECC",
X"E0C0",
X"DFC6",
X"E043",
X"DF49",
X"E0C0",
X"DAE4",
X"D8F0",
X"D873",
X"D873",
X"DC5B",
X"D6FC",
X"DAE4",
X"D7F6",
X"D508",
X"D67F",
X"D19D",
X"D96D",
X"D779",
X"D40E",
X"D6FC",
X"D96D",
X"DFC6",
X"E3AE",
X"E813",
X"EA84",
X"E98A",
X"EBFB",
X"ECF5",
X"EEE9",
X"F448",
X"F3CB",
X"F3CB",
X"F63C",
X"F34E",
X"F542",
X"F448",
X"F63C",
X"FB1E",
X"00FA",
X"036B",
X"0465",
X"06D6",
X"0659",
X"04E2",
X"0271",
X"FF06",
X"FD8F",
X"00FA",
X"02EE",
X"01F4",
X"007D",
X"FF06",
X"00FA",
X"FD8F",
X"FF06",
X"FF83",
X"FE89",
X"FD12",
X"FB1E",
X"FA24",
X"F9A7",
X"F63C",
X"F1D7",
X"F0DD",
X"F0DD",
X"EC78",
X"EF66",
X"EFE3",
X"EB01",
X"EDEF",
X"E90D",
X"E331",
X"E3AE",
X"E61F",
X"EA84",
X"EA07",
X"EA84",
X"EA07",
X"E61F",
X"E719",
X"E5A2",
X"E5A2",
X"E90D",
X"EC78",
X"EC78",
X"EE6C",
X"ED72",
X"ED72",
X"EDEF",
X"EDEF",
X"EF66",
X"F060",
X"F34E",
X"F254",
X"F0DD",
X"F4C5",
X"F6B9",
X"F8AD",
X"FF83",
X"03E8",
X"0947",
X"0A41",
X"0C35",
X"0C35",
X"0DAC",
X"0EA6",
X"1117",
X"1388",
X"14FF",
X"1B58",
X"1CCF",
X"186A",
X"15F9",
X"1964",
X"1D4C",
X"1D4C",
X"1FBD",
X"2134",
X"251C",
X"2B75",
X"2AF8",
X"2B75",
X"2EE0",
X"2BF2",
X"29FE",
X"2BF2",
X"324B",
X"32C8",
X"3633",
X"372D",
X"3633",
X"343F",
X"3151",
X"33C2",
X"2E63",
X"2D69",
X"30D4",
X"324B",
X"343F",
X"35B6",
X"324B",
X"31CE",
X"2CEC",
X"2B75",
X"2A7B",
X"2B75",
X"2E63",
X"2DE6",
X"2F5D",
X"2F5D",
X"2FDA",
X"2CEC",
X"2E63",
X"2D69",
X"2887",
X"251C",
X"249F",
X"1F40",
X"17ED",
X"101D",
X"0A41",
X"08CA",
X"01F4",
X"FD12",
X"FB9B",
X"FC95",
X"FC95",
X"F8AD",
X"F6B9",
X"F830",
X"F5BF",
X"F34E",
X"EFE3",
X"ED72",
X"E98A",
X"EA07",
X"E719",
X"DF49",
X"DA67",
X"D8F0",
X"DBDE",
X"E1BA",
X"E2B4",
X"E2B4",
X"E237",
X"DFC6",
X"DCD8",
X"DC5B",
X"DD55",
X"DC5B",
X"E043",
X"DFC6",
X"E1BA",
X"E237",
X"E4A8",
X"E90D",
X"EB7E",
X"EB7E",
X"EC78",
X"EA84",
X"F0DD",
X"F4C5",
X"F448",
X"F542",
X"F92A",
X"00FA",
X"04E2",
X"FC95",
X"00FA",
X"036B",
X"00FA",
X"05DC",
X"06D6",
X"07D0",
X"0947",
X"09C4",
X"0BB8",
X"0D2F",
X"101D",
X"0CB2",
X"0BB8",
X"0FA0",
X"0EA6",
X"0DAC",
X"101D",
X"1117",
X"0E29",
X"0ABE",
X"0ABE",
X"09C4",
X"084D",
X"0465",
X"FE89",
X"FD12",
X"FD8F",
X"FE89",
X"FE0C",
X"FB1E",
X"FA24",
X"FAA1",
X"F9A7",
X"F6B9",
X"F3CB",
X"F34E",
X"F254",
X"EFE3",
X"F1D7",
X"F15A",
X"F1D7",
X"EF66",
X"F254",
X"F448",
X"F34E",
X"F6B9",
X"F736",
X"F7B3",
X"F63C",
X"F5BF",
X"EF66",
X"F0DD",
X"EF66",
X"EA07",
X"E331",
X"DF49",
X"E2B4",
X"DF49",
X"DE4F",
X"DD55",
X"DE4F",
X"E61F",
X"E69C",
X"EDEF",
X"ECF5",
X"EA07",
X"E69C",
X"E3AE",
X"E2B4",
X"E890",
X"EB7E",
X"F060",
X"F2D1",
X"F5BF",
X"FA24",
X"FAA1",
X"F8AD",
X"FC95",
X"FD12",
X"FAA1",
X"FC95",
X"F9A7",
X"F92A",
X"F8AD",
X"F9A7",
X"FE89",
X"04E2",
X"05DC",
X"0659",
X"05DC",
X"055F",
X"0465",
X"FF83",
X"00FA",
X"0753",
X"0BB8",
X"109A",
X"1676",
X"14FF",
X"1388",
X"0CB2",
X"09C4",
X"0A41",
X"0A41",
X"0B3B",
X"101D",
X"0D2F",
X"0BB8",
X"0C35",
X"0A41",
X"055F",
X"07D0",
X"08CA",
X"084D",
X"03E8",
X"007D",
X"0177",
X"0465",
X"01F4",
X"05DC",
X"0B3B",
X"0ABE",
X"0EA6",
X"109A",
X"0E29",
X"101D",
X"0B3B",
X"084D",
X"06D6",
X"0A41",
X"0659",
X"055F",
X"0753",
X"07D0",
X"05DC",
X"02EE",
X"04E2",
X"05DC",
X"055F",
X"055F",
X"02EE",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"0177",
X"FC95",
X"FB9B",
X"FB1E",
X"FD8F",
X"FD12",
X"FD8F",
X"F9A7",
X"FA24",
X"F7B3",
X"F5BF",
X"F6B9",
X"F34E",
X"F63C",
X"F5BF",
X"F254",
X"F3CB",
X"F2D1",
X"F1D7",
X"EE6C",
X"EB01",
X"EB01",
X"EBFB",
X"EA84",
X"E813",
X"EC78",
X"EC78",
X"EB7E",
X"F0DD",
X"F254",
X"F34E",
X"F6B9",
X"F92A",
X"F9A7",
X"FE0C",
X"FF06",
X"00FA",
X"01F4",
X"03E8",
X"0271",
X"0177",
X"05DC",
X"0ABE",
X"09C4",
X"07D0",
X"0CB2",
X"1194",
X"1482",
X"15F9",
X"1482",
X"157C",
X"1964",
X"1A5E",
X"1DC9",
X"18E7",
X"186A",
X"17ED",
X"17ED",
X"18E7",
X"1CCF",
X"1B58",
X"1ADB",
X"1BD5",
X"17ED",
X"17ED",
X"128E",
X"1211",
X"1211",
X"109A",
X"0C35",
X"0B3B",
X"0CB2",
X"0A41",
X"08CA",
X"055F",
X"04E2",
X"04E2",
X"036B",
X"0271",
X"0271",
X"FD12",
X"01F4",
X"007D",
X"0271",
X"FC18",
X"FAA1",
X"0000",
X"FE89",
X"007D",
X"0271",
X"0271",
X"0271",
X"04E2",
X"055F",
X"03E8",
X"07D0",
X"07D0",
X"0753",
X"0465",
X"0177",
X"01F4",
X"02EE",
X"03E8",
X"036B",
X"0000",
X"0271",
X"04E2",
X"0271",
X"0271",
X"00FA",
X"02EE",
X"FE89",
X"0177",
X"0465",
X"0753",
X"06D6",
X"04E2",
X"0753",
X"03E8",
X"06D6",
X"0659",
X"0659",
X"036B",
X"01F4",
X"036B",
X"055F",
X"036B",
X"01F4",
X"0659",
X"055F",
X"036B",
X"05DC",
X"055F",
X"01F4",
X"FF06",
X"FD8F",
X"FC95",
X"FD12",
X"FD8F",
X"FA24",
X"F830",
X"F9A7",
X"F9A7",
X"F7B3",
X"F830",
X"F542",
X"EEE9",
X"EEE9",
X"F2D1",
X"F34E",
X"F15A",
X"EFE3",
X"F448",
X"F542",
X"F2D1",
X"F63C",
X"F736",
X"F7B3",
X"F6B9",
X"F448",
X"F5BF",
X"FB9B",
X"FC18",
X"FC95",
X"FAA1",
X"FF06",
X"FF06",
X"FC18",
X"FC95",
X"FF06",
X"FC18",
X"FE89",
X"FF83",
X"FD8F",
X"FA24",
X"FD8F",
X"FE0C",
X"FC18",
X"FB9B",
X"FB1E",
X"FE0C",
X"FAA1",
X"F542",
X"F3CB",
X"F448",
X"F5BF",
X"EFE3",
X"ED72",
X"EE6C",
X"EF66",
X"EEE9",
X"E719",
X"EA07",
X"E98A",
X"E69C",
X"E890",
X"E98A",
X"EA84",
X"EEE9",
X"ED72",
X"EBFB",
X"EDEF",
X"EDEF",
X"F060",
X"F2D1",
X"F2D1",
X"F254",
X"F448",
X"F2D1",
X"F736",
X"F5BF",
X"F63C",
X"F9A7",
X"FA24",
X"FB1E",
X"FB1E",
X"FC18",
X"F6B9",
X"F4C5",
X"FA24",
X"F6B9",
X"F63C",
X"F448",
X"FD12",
X"FD8F",
X"F9A7",
X"FF83",
X"036B",
X"055F",
X"03E8",
X"05DC",
X"01F4",
X"01F4",
X"055F",
X"0753",
X"055F",
X"05DC",
X"04E2",
X"0753",
X"01F4",
X"00FA",
X"FA24",
X"FA24",
X"FD12",
X"F63C",
X"F9A7",
X"FAA1",
X"FE89",
X"F92A",
X"FB1E",
X"FD8F",
X"FE0C",
X"FC18",
X"FE0C",
X"036B",
X"055F",
X"03E8",
X"03E8",
X"055F",
X"02EE",
X"FD12",
X"0271",
X"007D",
X"007D",
X"0271",
X"01F4",
X"0947",
X"036B",
X"07D0",
X"08CA",
X"0F23",
X"157C",
X"1405",
X"1211",
X"1388",
X"18E7",
X"18E7",
X"19E1",
X"1BD5",
X"1B58",
X"1676",
X"1DC9",
X"1EC3",
X"1964",
X"18E7",
X"186A",
X"1ADB",
X"18E7",
X"157C",
X"0EA6",
X"1482",
X"1194",
X"1388",
X"128E",
X"0A41",
X"0C35",
X"084D",
X"04E2",
X"04E2",
X"02EE",
X"0659",
X"0753",
X"05DC",
X"04E2",
X"0000",
X"FC18",
X"FB9B",
X"FB9B",
X"007D",
X"02EE",
X"FF06",
X"02EE",
X"007D",
X"01F4",
X"FE0C",
X"FF06",
X"03E8",
X"FE89",
X"FF83",
X"0177",
X"FF06",
X"FD12",
X"FB1E",
X"FAA1",
X"FD8F",
X"FB1E",
X"FA24",
X"FE0C",
X"FC18",
X"FE0C",
X"FE0C",
X"FE0C",
X"01F4",
X"01F4",
X"0271",
X"01F4",
X"0177",
X"0177",
X"03E8",
X"0271",
X"0271",
X"0659",
X"055F",
X"036B",
X"007D",
X"00FA",
X"FC95",
X"F9A7",
X"F7B3",
X"F7B3",
X"F9A7",
X"00FA",
X"0000",
X"FD8F",
X"FF06",
X"FAA1",
X"FAA1",
X"FD8F",
X"F9A7",
X"FC18",
X"F9A7",
X"F8AD",
X"FD12",
X"F830",
X"FB1E",
X"FA24",
X"F736",
X"FB1E",
X"FE89",
X"F8AD",
X"F830",
X"F736",
X"F6B9",
X"FC18",
X"FC18",
X"F9A7",
X"FE0C",
X"FE89",
X"FE0C",
X"FE89",
X"0177",
X"0465",
X"05DC",
X"055F",
X"055F",
X"0947",
X"0B3B",
X"07D0",
X"07D0",
X"09C4",
X"0BB8",
X"0B3B",
X"08CA",
X"0753",
X"08CA",
X"09C4",
X"0B3B",
X"0B3B",
X"0CB2",
X"0E29",
X"0C35",
X"0E29",
X"0A41",
X"08CA",
X"04E2",
X"055F",
X"05DC",
X"055F",
X"06D6",
X"02EE",
X"01F4",
X"036B",
X"0177",
X"02EE",
X"FE89",
X"02EE",
X"007D",
X"0000",
X"04E2",
X"03E8",
X"04E2",
X"036B",
X"01F4",
X"0000",
X"03E8",
X"FE0C",
X"036B",
X"06D6",
X"01F4",
X"036B",
X"036B",
X"0465",
X"0947",
X"0A41",
X"0F23",
X"1117",
X"1405",
X"0DAC",
X"0CB2",
X"0CB2",
X"0C35",
X"0947",
X"0C35",
X"0659",
X"05DC",
X"07D0",
X"0C35",
X"0947",
X"0A41",
X"0E29",
X"0E29",
X"0C35",
X"09C4",
X"0DAC",
X"0D2F",
X"09C4",
X"09C4",
X"0D2F",
X"02EE",
X"FB1E",
X"F9A7",
X"F5BF",
X"F254",
X"F6B9",
X"EDEF",
X"EDEF",
X"EB01",
X"EA07",
X"EBFB",
X"EA84",
X"E61F",
X"E5A2",
X"E796",
X"E69C",
X"E237",
X"E043",
X"E4A8",
X"E719",
X"E890",
X"E90D",
X"E69C",
X"E525",
X"E98A",
X"E719",
X"E98A",
X"EB7E",
X"EBFB",
X"EDEF",
X"EB7E",
X"EA84",
X"EA07",
X"EE6C",
X"F2D1",
X"F4C5",
X"F448",
X"F542",
X"F3CB",
X"F3CB",
X"F542",
X"F7B3",
X"F830",
X"F92A",
X"F7B3",
X"FAA1",
X"FD12",
X"FB9B",
X"FC95",
X"FB1E",
X"F8AD",
X"F92A",
X"F736",
X"F7B3",
X"F448",
X"F4C5",
X"F254",
X"F1D7",
X"F2D1",
X"F254",
X"F0DD",
X"ECF5",
X"F15A",
X"F060",
X"F254",
X"F0DD",
X"F1D7",
X"ECF5",
X"EEE9",
X"F3CB",
X"F1D7",
X"EFE3",
X"F0DD",
X"F2D1",
X"F542",
X"F5BF",
X"F4C5",
X"F3CB",
X"F448",
X"F5BF",
X"F5BF",
X"F542",
X"F3CB",
X"F448",
X"F3CB",
X"F63C",
X"F15A",
X"F15A",
X"F4C5",
X"F542",
X"F34E",
X"F34E",
X"F1D7",
X"F254",
X"F2D1",
X"F542",
X"F63C",
X"F34E",
X"F448",
X"F3CB",
X"F3CB",
X"F542",
X"F63C",
X"F3CB",
X"F34E",
X"F254",
X"F1D7",
X"F15A",
X"F34E",
X"F542",
X"F830",
X"F92A",
X"F8AD",
X"F9A7",
X"FB9B",
X"FC95",
X"FC95",
X"FC18",
X"FF06",
X"01F4",
X"00FA",
X"036B",
X"055F",
X"08CA",
X"0A41",
X"0BB8",
X"0F23",
X"1194",
X"1194",
X"1388",
X"157C",
X"17ED",
X"1B58",
X"1BD5",
X"1D4C",
X"1D4C",
X"1BD5",
X"1CCF",
X"2134",
X"2599",
X"251C",
X"2693",
X"2981",
X"278D",
X"2710",
X"2981",
X"2BF2",
X"29FE",
X"2887",
X"2981",
X"29FE",
X"2C6F",
X"2904",
X"2422",
X"2710",
X"2710",
X"280A",
X"23A5",
X"1F40",
X"20B7",
X"1E46",
X"1DC9",
X"1CCF",
X"1964",
X"17ED",
X"186A",
X"1770",
X"1770",
X"1676",
X"157C",
X"186A",
X"16F3",
X"1405",
X"128E",
X"109A",
X"0ABE",
X"084D",
X"08CA",
X"08CA",
X"04E2",
X"02EE",
X"0465",
X"02EE",
X"007D",
X"0271",
X"02EE",
X"02EE",
X"0271",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"0271",
X"0000",
X"0271",
X"00FA",
X"0177",
X"00FA",
X"FE0C",
X"FC95",
X"FE89",
X"FF06",
X"FE89",
X"007D",
X"01F4",
X"055F",
X"084D",
X"0BB8",
X"084D",
X"0659",
X"0D2F",
X"09C4",
X"0947",
X"055F",
X"0753",
X"084D",
X"0659",
X"0659",
X"055F",
X"0ABE",
X"09C4",
X"09C4",
X"0CB2",
X"0D2F",
X"0B3B",
X"0C35",
X"0D2F",
X"0CB2",
X"0BB8",
X"0DAC",
X"0C35",
X"09C4",
X"0BB8",
X"09C4",
X"04E2",
X"03E8",
X"04E2",
X"0465",
X"06D6",
X"036B",
X"007D",
X"FC18",
X"FD12",
X"FAA1",
X"FB9B",
X"F92A",
X"F4C5",
X"F3CB",
X"F542",
X"F3CB",
X"F4C5",
X"F4C5",
X"F2D1",
X"F060",
X"ECF5",
X"EB7E",
X"EF66",
X"F15A",
X"F0DD",
X"ECF5",
X"F060",
X"EC78",
X"EBFB",
X"EEE9",
X"E90D",
X"E890",
X"E61F",
X"E3AE",
X"E331",
X"DFC6",
X"DECC",
X"DE4F",
X"DDD2",
X"DE4F",
X"D96D",
X"DAE4",
X"DC5B",
X"DDD2",
X"DB61",
X"DA67",
X"DA67",
X"D9EA",
X"DB61",
X"D7F6",
X"D67F",
X"DA67",
X"D602",
X"DAE4",
X"D9EA",
X"DA67",
X"E043",
X"DB61",
X"DECC",
X"DB61",
X"DAE4",
X"DECC",
X"DE4F",
X"E0C0",
X"E0C0",
X"DE4F",
X"E0C0",
X"E1BA",
X"DFC6",
X"E525",
X"E42B",
X"E4A8",
X"E3AE",
X"E4A8",
X"E61F",
X"E890",
X"ED72",
X"EEE9",
X"F15A",
X"F34E",
X"F34E",
X"F4C5",
X"F9A7",
X"FB1E",
X"FA24",
X"FC95",
X"FC95",
X"FC18",
X"FE89",
X"FB9B",
X"FAA1",
X"FF06",
X"01F4",
X"04E2",
X"0B3B",
X"09C4",
X"0ABE",
X"0D2F",
X"0B3B",
X"0D2F",
X"0B3B",
X"0B3B",
X"0EA6",
X"0E29",
X"1194",
X"1194",
X"1117",
X"15F9",
X"130B",
X"101D",
X"0EA6",
X"0F23",
X"128E",
X"128E",
X"1211",
X"1482",
X"1405",
X"128E",
X"1211",
X"0F23",
X"1194",
X"1194",
X"0F23",
X"101D",
X"0F23",
X"0F23",
X"128E",
X"0EA6",
X"1405",
X"128E",
X"1117",
X"157C",
X"1405",
X"1482",
X"14FF",
X"1388",
X"14FF",
X"15F9",
X"1405",
X"157C",
X"1405",
X"1117",
X"1482",
X"1482",
X"15F9",
X"128E",
X"109A",
X"128E",
X"0F23",
X"109A",
X"109A",
X"1211",
X"14FF",
X"1676",
X"14FF",
X"1482",
X"128E",
X"157C",
X"15F9",
X"1405",
X"130B",
X"128E",
X"1388",
X"128E",
X"101D",
X"128E",
X"1388",
X"1117",
X"1388",
X"1211",
X"0E29",
X"0C35",
X"0B3B",
X"0C35",
X"0C35",
X"09C4",
X"0947",
X"0A41",
X"0753",
X"0659",
X"084D",
X"01F4",
X"FF06",
X"007D",
X"0000",
X"FD12",
X"FF06",
X"FC95",
X"FB1E",
X"F92A",
X"F736",
X"F830",
X"F830",
X"F736",
X"F6B9",
X"F4C5",
X"F2D1",
X"F2D1",
X"F0DD",
X"F060",
X"EE6C",
X"EFE3",
X"F15A",
X"EF66",
X"ECF5",
X"EFE3",
X"EE6C",
X"EBFB",
X"EBFB",
X"EEE9",
X"ED72",
X"EBFB",
X"EE6C",
X"F34E",
X"F63C",
X"F6B9",
X"F9A7",
X"F736",
X"F63C",
X"F9A7",
X"FC95",
X"FC18",
X"F8AD",
X"F9A7",
X"FC18",
X"FD12",
X"FC95",
X"FC95",
X"FA24",
X"F8AD",
X"F92A",
X"F6B9",
X"F92A",
X"F830",
X"FAA1",
X"FC95",
X"FB9B",
X"FE89",
X"007D",
X"00FA",
X"00FA",
X"0000",
X"0271",
X"00FA",
X"01F4",
X"04E2",
X"0465",
X"01F4",
X"03E8",
X"05DC",
X"06D6",
X"0465",
X"0465",
X"03E8",
X"0465",
X"07D0",
X"05DC",
X"0465",
X"03E8",
X"06D6",
X"07D0",
X"08CA",
X"06D6",
X"0947",
X"09C4",
X"0ABE",
X"08CA",
X"05DC",
X"0753",
X"084D",
X"03E8",
X"0177",
X"01F4",
X"007D",
X"00FA",
X"00FA",
X"0271",
X"0177",
X"036B",
X"036B",
X"03E8",
X"036B",
X"0271",
X"0271",
X"0271",
X"FE0C",
X"FE89",
X"FD8F",
X"FC95",
X"FC95",
X"F9A7",
X"F6B9",
X"F3CB",
X"F92A",
X"F15A",
X"EDEF",
X"F542",
X"F830",
X"F448",
X"EB01",
X"F2D1",
X"F448",
X"EEE9",
X"F15A",
X"F34E",
X"EE6C",
X"E98A",
X"EE6C",
X"F2D1",
X"EDEF",
X"EB7E",
X"EEE9",
X"ED72",
X"ECF5",
X"EE6C",
X"EE6C",
X"EB01",
X"EA07",
X"EDEF",
X"ECF5",
X"EB7E",
X"EBFB",
X"EBFB",
X"F0DD",
X"F2D1",
X"EE6C",
X"F1D7",
X"F34E",
X"F34E",
X"FA24",
X"F6B9",
X"F5BF",
X"FC95",
X"FD8F",
X"FD8F",
X"FC18",
X"FF06",
X"007D",
X"02EE",
X"05DC",
X"09C4",
X"0947",
X"09C4",
X"0CB2",
X"101D",
X"1482",
X"128E",
X"101D",
X"1117",
X"14FF",
X"16F3",
X"16F3",
X"19E1",
X"1BD5",
X"1C52",
X"1BD5",
X"1DC9",
X"1F40",
X"20B7",
X"203A",
X"20B7",
X"203A",
X"1E46",
X"1D4C",
X"1B58",
X"1BD5",
X"1A5E",
X"186A",
X"1676",
X"14FF",
X"1482",
X"1194",
X"1211",
X"101D",
X"0C35",
X"0A41",
X"0B3B",
X"0E29",
X"0947",
X"036B",
X"036B",
X"02EE",
X"036B",
X"FE89",
X"FAA1",
X"FA24",
X"F7B3",
X"F830",
X"FC95",
X"FB9B",
X"FA24",
X"F8AD",
X"F8AD",
X"F92A",
X"F9A7",
X"F9A7",
X"F8AD",
X"F92A",
X"FA24",
X"F8AD",
X"F6B9",
X"F7B3",
X"F8AD",
X"F6B9",
X"F8AD",
X"F8AD",
X"F92A",
X"F92A",
X"FAA1",
X"FB9B",
X"FB1E",
X"FB9B",
X"FD12",
X"0271",
X"0271",
X"04E2",
X"055F",
X"0465",
X"05DC",
X"0947",
X"0A41",
X"0ABE",
X"0A41",
X"0ABE",
X"0A41",
X"09C4",
X"06D6",
X"0753",
X"07D0",
X"04E2",
X"0271",
X"0271",
X"00FA",
X"FC18",
X"FF06",
X"FE0C",
X"FC18",
X"FC18",
X"FD8F",
X"FE0C",
X"F9A7",
X"F92A",
X"F8AD",
X"F542",
X"F63C",
X"F542",
X"F448",
X"F2D1",
X"F1D7",
X"F34E",
X"F060",
X"EDEF",
X"EBFB",
X"EBFB",
X"EE6C",
X"EA84",
X"E98A",
X"EF66",
X"E890",
X"EA07",
X"EBFB",
X"EDEF",
X"EFE3",
X"ECF5",
X"F4C5",
X"F3CB",
X"F254",
X"F1D7",
X"F15A",
X"F542",
X"F7B3",
X"F542",
X"F4C5",
X"F92A",
X"FC18",
X"FAA1",
X"F92A",
X"F9A7",
X"FC95",
X"FE0C",
X"FC95",
X"FD12",
X"FB9B",
X"FE89",
X"FC18",
X"FE89",
X"0177",
X"FD12",
X"FC95",
X"FF83",
X"FE0C",
X"F92A",
X"F92A",
X"FAA1",
X"F9A7",
X"FB1E",
X"FD12",
X"FC95",
X"FC18",
X"FC95",
X"FD8F",
X"FC95",
X"FD12",
X"F92A",
X"F8AD",
X"F7B3",
X"F542",
X"F4C5",
X"F542",
X"F542",
X"F1D7",
X"F060",
X"F2D1",
X"F2D1",
X"EFE3",
X"F15A",
X"F060",
X"F0DD",
X"F34E",
X"F34E",
X"F4C5",
X"F448",
X"F254",
X"F34E",
X"F448",
X"FA24",
X"F8AD",
X"F736",
X"FAA1",
X"FC95",
X"FE89",
X"FC95",
X"FF06",
X"007D",
X"FF83",
X"0000",
X"036B",
X"0659",
X"0753",
X"0B3B",
X"0C35",
X"1211",
X"1482",
X"1676",
X"1ADB",
X"1E46",
X"1E46",
X"1C52",
X"1EC3",
X"1C52",
X"1BD5",
X"1CCF",
X"1EC3",
X"21B1",
X"222E",
X"2328",
X"222E",
X"2599",
X"2710",
X"2693",
X"278D",
X"2981",
X"2887",
X"2710",
X"2616",
X"2693",
X"2616",
X"2693",
X"2422",
X"203A",
X"1DC9",
X"1D4C",
X"17ED",
X"1211",
X"128E",
X"0D2F",
X"0BB8",
X"084D",
X"055F",
X"02EE",
X"FE89",
X"0000",
X"FE89",
X"FB9B",
X"F736",
X"FC95",
X"FB9B",
X"F63C",
X"FB1E",
X"FAA1",
X"F92A",
X"F3CB",
X"F6B9",
X"F3CB",
X"ED72",
X"EEE9",
X"EF66",
X"ECF5",
X"EB01",
X"EBFB",
X"ECF5",
X"ED72",
X"ECF5",
X"EBFB",
X"ECF5",
X"EF66",
X"F060",
X"F448",
X"F254",
X"F2D1",
X"F542",
X"F2D1",
X"F4C5",
X"F8AD",
X"F5BF",
X"F92A",
X"FD12",
X"00FA",
X"007D",
X"FE89",
X"01F4",
X"007D",
X"FE0C",
X"FF06",
X"FF06",
X"FF83",
X"FF06",
X"FD8F",
X"FD12",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"FD8F",
X"007D",
X"00FA",
X"0000",
X"0177",
X"FF83",
X"0000",
X"FF83",
X"0271",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FC95",
X"FB9B",
X"FB9B",
X"F9A7",
X"F92A",
X"F6B9",
X"F254",
X"F15A",
X"F254",
X"EF66",
X"F060",
X"F060",
X"EDEF",
X"EE6C",
X"EE6C",
X"EEE9",
X"EFE3",
X"F542",
X"F060",
X"ED72",
X"F736",
X"EF66",
X"EFE3",
X"F15A",
X"ED72",
X"F34E",
X"F1D7",
X"EBFB",
X"F1D7",
X"F0DD",
X"F060",
X"F448",
X"F7B3",
X"F92A",
X"F92A",
X"FD8F",
X"FD8F",
X"FF06",
X"FE89",
X"02EE",
X"06D6",
X"036B",
X"0659",
X"09C4",
X"08CA",
X"0947",
X"0D2F",
X"109A",
X"101D",
X"1211",
X"1211",
X"1482",
X"1676",
X"1676",
X"1770",
X"1770",
X"157C",
X"17ED",
X"186A",
X"1676",
X"14FF",
X"157C",
X"1676",
X"1211",
X"0D2F",
X"0EA6",
X"0DAC",
X"0BB8",
X"0EA6",
X"0CB2",
X"0BB8",
X"0ABE",
X"0947",
X"07D0",
X"04E2",
X"05DC",
X"06D6",
X"03E8",
X"01F4",
X"FF83",
X"FD12",
X"FB9B",
X"FB1E",
X"FB9B",
X"FAA1",
X"F9A7",
X"F8AD",
X"F6B9",
X"F8AD",
X"F7B3",
X"F6B9",
X"F5BF",
X"F830",
X"F7B3",
X"F92A",
X"FB1E",
X"F7B3",
X"FF83",
X"FE0C",
X"FAA1",
X"01F4",
X"FF06",
X"0177",
X"FE0C",
X"FF06",
X"0177",
X"FD8F",
X"01F4",
X"0000",
X"FF06",
X"055F",
X"0465",
X"00FA",
X"03E8",
X"02EE",
X"04E2",
X"0659",
X"03E8",
X"007D",
X"0271",
X"01F4",
X"0271",
X"FE0C",
X"FE89",
X"FD8F",
X"F92A",
X"FF06",
X"F542",
X"FAA1",
X"F830",
X"F4C5",
X"F5BF",
X"EFE3",
X"F34E",
X"F254",
X"EF66",
X"ECF5",
X"EDEF",
X"EFE3",
X"EEE9",
X"EF66",
X"F0DD",
X"F15A",
X"F0DD",
X"F1D7",
X"F060",
X"EE6C",
X"EFE3",
X"EEE9",
X"ED72",
X"ECF5",
X"F060",
X"EF66",
X"EC78",
X"EEE9",
X"EE6C",
X"EFE3",
X"EFE3",
X"F254",
X"F1D7",
X"F5BF",
X"F6B9",
X"F5BF",
X"F5BF",
X"F7B3",
X"F6B9",
X"F5BF",
X"F63C",
X"F542",
X"F6B9",
X"F92A",
X"FC18",
X"FD12",
X"FE89",
X"02EE",
X"0177",
X"00FA",
X"0177",
X"0177",
X"01F4",
X"007D",
X"FE89",
X"FD8F",
X"FD12",
X"FA24",
X"FB9B",
X"F92A",
X"F92A",
X"FAA1",
X"FF06",
X"007D",
X"0000",
X"007D",
X"02EE",
X"01F4",
X"02EE",
X"036B",
X"01F4",
X"036B",
X"036B",
X"02EE",
X"0659",
X"06D6",
X"07D0",
X"08CA",
X"084D",
X"08CA",
X"05DC",
X"0659",
X"04E2",
X"036B",
X"06D6",
X"0465",
X"08CA",
X"0A41",
X"0659",
X"08CA",
X"0C35",
X"0ABE",
X"0ABE",
X"0DAC",
X"0BB8",
X"0F23",
X"0F23",
X"0FA0",
X"0EA6",
X"0D2F",
X"0EA6",
X"0CB2",
X"0D2F",
X"0FA0",
X"0D2F",
X"101D",
X"0F23",
X"0F23",
X"0D2F",
X"109A",
X"0DAC",
X"0C35",
X"0DAC",
X"0DAC",
X"0F23",
X"0EA6",
X"1194",
X"128E",
X"1194",
X"101D",
X"128E",
X"1211",
X"1117",
X"128E",
X"1482",
X"14FF",
X"130B",
X"1388",
X"130B",
X"157C",
X"14FF",
X"14FF",
X"15F9",
X"1676",
X"15F9",
X"1388",
X"157C",
X"18E7",
X"186A",
X"186A",
X"1964",
X"1770",
X"15F9",
X"1482",
X"16F3",
X"1482",
X"1405",
X"128E",
X"1211",
X"109A",
X"0D2F",
X"0CB2",
X"0A41",
X"07D0",
X"07D0",
X"04E2",
X"0465",
X"02EE",
X"0177",
X"0271",
X"02EE",
X"0177",
X"007D",
X"01F4",
X"007D",
X"0000",
X"FF83",
X"0000",
X"0000",
X"0000",
X"FC95",
X"FB9B",
X"FB1E",
X"F92A",
X"F9A7",
X"FB1E",
X"F9A7",
X"FB9B",
X"FD12",
X"0000",
X"0000",
X"0000",
X"FE89",
X"FD12",
X"FD12",
X"FB1E",
X"FA24",
X"F8AD",
X"F736",
X"F63C",
X"F7B3",
X"F830",
X"F7B3",
X"F7B3",
X"F830",
X"F63C",
X"F542",
X"F6B9",
X"F6B9",
X"F448",
X"F4C5",
X"F2D1",
X"F3CB",
X"F34E",
X"F254",
X"F15A",
X"EE6C",
X"EEE9",
X"ED72",
X"EB7E",
X"EE6C",
X"EC78",
X"EA07",
X"EBFB",
X"E98A",
X"EB7E",
X"EBFB",
X"E90D",
X"E98A",
X"EA07",
X"E98A",
X"EA84",
X"E813",
X"E719",
X"E69C",
X"E42B",
X"E42B",
X"E331",
X"E237",
X"E237",
X"E2B4",
X"E331",
X"E42B",
X"E525",
X"E42B",
X"E61F",
X"E69C",
X"E719",
X"E890",
X"E813",
X"E61F",
X"E5A2",
X"E69C",
X"E525",
X"E61F",
X"E69C",
X"E719",
X"EA84",
X"EA07",
X"EB01",
X"EB7E",
X"EB01",
X"EBFB",
X"EB7E",
X"EB7E",
X"EA07",
X"EA07",
X"EC78",
X"EC78",
X"EBFB",
X"EE6C",
X"EC78",
X"EFE3",
X"EEE9",
X"EE6C",
X"F254",
X"F060",
X"F254",
X"F448",
X"F448",
X"F6B9",
X"F736",
X"F92A",
X"FA24",
X"FB1E",
X"FB9B",
X"FB1E",
X"FAA1",
X"FA24",
X"FAA1",
X"F8AD",
X"F8AD",
X"F830",
X"F92A",
X"F92A",
X"F92A",
X"FD8F",
X"FE89",
X"FD12",
X"FE0C",
X"007D",
X"00FA",
X"036B",
X"04E2",
X"055F",
X"05DC",
X"0947",
X"09C4",
X"0C35",
X"0BB8",
X"084D",
X"09C4",
X"0DAC",
X"0D2F",
X"0BB8",
X"0C35",
X"0C35",
X"0DAC",
X"0DAC",
X"0EA6",
X"1388",
X"15F9",
X"15F9",
X"16F3",
X"1C52",
X"1DC9",
X"1DC9",
X"22AB",
X"2328",
X"2134",
X"222E",
X"22AB",
X"2422",
X"23A5",
X"249F",
X"2599",
X"22AB",
X"22AB",
X"2328",
X"2599",
X"2887",
X"251C",
X"2599",
X"2904",
X"2887",
X"278D",
X"2981",
X"2B75",
X"29FE",
X"2887",
X"2C6F",
X"2D69",
X"29FE",
X"249F",
X"2616",
X"280A",
X"23A5",
X"21B1",
X"22AB",
X"222E",
X"1F40",
X"1EC3",
X"1DC9",
X"1ADB",
X"1770",
X"157C",
X"130B",
X"1117",
X"109A",
X"1211",
X"128E",
X"0E29",
X"0C35",
X"0D2F",
X"0C35",
X"0ABE",
X"0753",
X"05DC",
X"08CA",
X"0659",
X"03E8",
X"05DC",
X"02EE",
X"FF83",
X"0177",
X"FF83",
X"FC18",
X"FC18",
X"0000",
X"01F4",
X"FE89",
X"007D",
X"FE0C",
X"FE0C",
X"FF06",
X"FE0C",
X"FB9B",
X"FA24",
X"FA24",
X"F8AD",
X"F92A",
X"F92A",
X"FB1E",
X"FA24",
X"FF06",
X"0000",
X"FB9B",
X"FE89",
X"FC95",
X"F8AD",
X"FC95",
X"FAA1",
X"FAA1",
X"F92A",
X"F736",
X"F92A",
X"F7B3",
X"F542",
X"F4C5",
X"F3CB",
X"F060",
X"EEE9",
X"EB7E",
X"EBFB",
X"ECF5",
X"EA84",
X"EB7E",
X"ECF5",
X"ED72",
X"E890",
X"E525",
X"E719",
X"E5A2",
X"E719",
X"E5A2",
X"E69C",
X"E42B",
X"E3AE",
X"E331",
X"E5A2",
X"E796",
X"E3AE",
X"E5A2",
X"E813",
X"E98A",
X"E719",
X"E813",
X"E98A",
X"E98A",
X"EA84",
X"EBFB",
X"EA84",
X"EB7E",
X"EC78",
X"ECF5",
X"EE6C",
X"EE6C",
X"EE6C",
X"EDEF",
X"F15A",
X"F0DD",
X"F1D7",
X"F254",
X"F1D7",
X"F1D7",
X"F34E",
X"F2D1",
X"F15A",
X"F1D7",
X"F15A",
X"F15A",
X"F1D7",
X"F448",
X"F254",
X"F1D7",
X"F15A",
X"F3CB",
X"F0DD",
X"F060",
X"F2D1",
X"F1D7",
X"F15A",
X"F0DD",
X"F0DD",
X"F0DD",
X"EF66",
X"EF66",
X"EC78",
X"ECF5",
X"ECF5",
X"EB7E",
X"EDEF",
X"EDEF",
X"EF66",
X"EDEF",
X"EEE9",
X"EDEF",
X"EE6C",
X"F060",
X"F060",
X"EFE3",
X"EF66",
X"F15A",
X"F060",
X"F0DD",
X"F448",
X"F34E",
X"F0DD",
X"F34E",
X"F5BF",
X"F3CB",
X"F542",
X"F542",
X"F63C",
X"F7B3",
X"FC18",
X"FC18",
X"FD12",
X"0000",
X"FF83",
X"00FA",
X"0271",
X"02EE",
X"0271",
X"055F",
X"06D6",
X"0753",
X"0947",
X"0ABE",
X"0FA0",
X"0EA6",
X"1117",
X"15F9",
X"1211",
X"1405",
X"14FF",
X"16F3",
X"157C",
X"1676",
X"18E7",
X"19E1",
X"1B58",
X"1ADB",
X"19E1",
X"1A5E",
X"1DC9",
X"1D4C",
X"1CCF",
X"1E46",
X"1D4C",
X"1D4C",
X"1F40",
X"1F40",
X"1E46",
X"1DC9",
X"1B58",
X"1964",
X"18E7",
X"1964",
X"1770",
X"15F9",
X"17ED",
X"14FF",
X"14FF",
X"17ED",
X"17ED",
X"157C",
X"1405",
X"128E",
X"1117",
X"1117",
X"109A",
X"101D",
X"0F23",
X"0FA0",
X"0F23",
X"0F23",
X"0E29",
X"0F23",
X"109A",
X"0FA0",
X"0FA0",
X"128E",
X"109A",
X"0FA0",
X"101D",
X"101D",
X"1211",
X"109A",
X"1117",
X"109A",
X"1194",
X"109A",
X"1194",
X"1388",
X"1482",
X"15F9",
X"15F9",
X"15F9",
X"157C",
X"1388",
X"1211",
X"1211",
X"130B",
X"1194",
X"0FA0",
X"0FA0",
X"0FA0",
X"0E29",
X"0EA6",
X"0C35",
X"0ABE",
X"0A41",
X"0947",
X"05DC",
X"0753",
X"04E2",
X"055F",
X"02EE",
X"036B",
X"0753",
X"02EE",
X"05DC",
X"05DC",
X"0271",
X"04E2",
X"03E8",
X"02EE",
X"036B",
X"0271",
X"036B",
X"0000",
X"FF06",
X"007D",
X"FF06",
X"FF06",
X"FB1E",
X"FAA1",
X"F8AD",
X"F9A7",
X"F63C",
X"F63C",
X"F4C5",
X"F34E",
X"EF66",
X"F736",
X"F254",
X"EA07",
X"F060",
X"F15A",
X"EC78",
X"E813",
X"ED72",
X"EC78",
X"E90D",
X"E719",
X"E69C",
X"E4A8",
X"E890",
X"E237",
X"DD55",
X"E61F",
X"DECC",
X"DECC",
X"DECC",
X"DBDE",
X"E4A8",
X"DAE4",
X"DE4F",
X"E0C0",
X"DCD8",
X"E237",
X"E0C0",
X"DFC6",
X"E043",
X"DF49",
X"DFC6",
X"DD55",
X"DECC",
X"DE4F",
X"DECC",
X"DFC6",
X"E0C0",
X"E043",
X"E1BA",
X"E3AE",
X"E237",
X"E331",
X"E525",
X"E4A8",
X"E525",
X"E525",
X"E4A8",
X"E61F",
X"E796",
X"EA07",
X"EA07",
X"EC78",
X"EEE9",
X"EDEF",
X"EEE9",
X"EFE3",
X"F0DD",
X"F15A",
X"F1D7",
X"F448",
X"F448",
X"F34E",
X"F4C5",
X"F254",
X"F3CB",
X"F6B9",
X"F7B3",
X"F736",
X"F830",
X"FB9B",
X"FC18",
X"FB1E",
X"FC95",
X"FE89",
X"FD8F",
X"0271",
X"01F4",
X"0271",
X"0271",
X"036B",
X"0465",
X"02EE",
X"01F4",
X"036B",
X"04E2",
X"055F",
X"0659",
X"09C4",
X"0BB8",
X"0ABE",
X"0B3B",
X"0CB2",
X"0DAC",
X"0C35",
X"0CB2",
X"0E29",
X"0BB8",
X"0ABE",
X"0A41",
X"0A41",
X"07D0",
X"0947",
X"0ABE",
X"0A41",
X"0947",
X"0A41",
X"0B3B",
X"0CB2",
X"0B3B",
X"0ABE",
X"0B3B",
X"0D2F",
X"0D2F",
X"0E29",
X"0EA6",
X"0EA6",
X"1194",
X"101D",
X"0FA0",
X"1117",
X"109A",
X"0EA6",
X"1211",
X"0F23",
X"1117",
X"130B",
X"1117",
X"128E",
X"130B",
X"15F9",
X"1770",
X"18E7",
X"16F3",
X"186A",
X"1964",
X"1A5E",
X"1A5E",
X"1ADB",
X"1B58",
X"1CCF",
X"1C52",
X"1D4C",
X"1E46",
X"1EC3",
X"203A",
X"2134",
X"1FBD",
X"203A",
X"22AB",
X"20B7",
X"1FBD",
X"20B7",
X"2134",
X"1DC9",
X"1D4C",
X"1F40",
X"1FBD",
X"1F40",
X"1EC3",
X"1FBD",
X"1E46",
X"1CCF",
X"1BD5",
X"19E1",
X"1964",
X"1770",
X"1388",
X"1388",
X"1117",
X"0FA0",
X"0DAC",
X"0E29",
X"0D2F",
X"0CB2",
X"0BB8",
X"0B3B",
X"0B3B",
X"0A41",
X"0947",
X"0753",
X"06D6",
X"055F",
X"0271",
X"01F4",
X"00FA",
X"FE0C",
X"FC18",
X"FC18",
X"F92A",
X"F9A7",
X"FC18",
X"FAA1",
X"F92A",
X"FC95",
X"FB1E",
X"FB1E",
X"FB1E",
X"FAA1",
X"F736",
X"F92A",
X"F8AD",
X"F6B9",
X"F5BF",
X"F0DD",
X"F34E",
X"F0DD",
X"EF66",
X"EDEF",
X"ED72",
X"EFE3",
X"ED72",
X"EA84",
X"EA84",
X"EA07",
X"E90D",
X"E5A2",
X"E69C",
X"E5A2",
X"E525",
X"DF49",
X"E2B4",
X"DDD2",
X"DCD8",
X"DD55",
X"D602",
X"E0C0",
X"D873",
X"D314",
X"DBDE",
X"DE4F",
X"DB61",
X"D7F6",
X"D585",
X"D779",
X"DF49",
X"E043",
X"DBDE",
X"D6FC",
X"E043",
X"DC5B",
X"DE4F",
X"E331",
X"E1BA",
X"DFC6",
X"DBDE",
X"E42B",
X"E813",
X"E0C0",
X"E5A2",
X"EDEF",
X"EA07",
X"EBFB",
X"E61F",
X"EB7E",
X"F060",
X"F1D7",
X"F2D1",
X"F254",
X"F8AD",
X"F4C5",
X"F448",
X"F9A7",
X"FB9B",
X"FB1E",
X"FC95",
X"FE89",
X"FF06",
X"03E8",
X"0659",
X"02EE",
X"05DC",
X"0753",
X"0BB8",
X"0BB8",
X"0A41",
X"0ABE",
X"0CB2",
X"0B3B",
X"0ABE",
X"09C4",
X"0A41",
X"09C4",
X"07D0",
X"0753",
X"0947",
X"09C4",
X"0753",
X"07D0",
X"0659",
X"06D6",
X"0753",
X"05DC",
X"0659",
X"0753",
X"0659",
X"05DC",
X"03E8",
X"01F4",
X"007D",
X"0000",
X"FD8F",
X"FC95",
X"FB1E",
X"F9A7",
X"F92A",
X"F92A",
X"F9A7",
X"FA24",
X"FC18",
X"F8AD",
X"F830",
X"FC95",
X"FF06",
X"FF83",
X"FB9B",
X"0000",
X"FF83",
X"0000",
X"01F4",
X"01F4",
X"FF06",
X"FF83",
X"04E2",
X"007D",
X"FE89",
X"00FA",
X"0465",
X"06D6",
X"055F",
X"0753",
X"06D6",
X"08CA",
X"0BB8",
X"0B3B",
X"0CB2",
X"0ABE",
X"09C4",
X"0DAC",
X"1117",
X"1211",
X"128E",
X"1194",
X"130B",
X"1388",
X"1211",
X"1211",
X"1194",
X"1388",
X"1211",
X"1405",
X"1211",
X"1194",
X"0F23",
X"0FA0",
X"1482",
X"128E",
X"1211",
X"130B",
X"1388",
X"1405",
X"15F9",
X"1194",
X"0F23",
X"130B",
X"14FF",
X"157C",
X"128E",
X"101D",
X"101D",
X"1194",
X"101D",
X"0F23",
X"0EA6",
X"0EA6",
X"0F23",
X"101D",
X"0EA6",
X"0FA0",
X"128E",
X"128E",
X"101D",
X"101D",
X"1211",
X"1388",
X"1388",
X"130B",
X"1194",
X"101D",
X"1388",
X"1211",
X"1388",
X"1117",
X"0E29",
X"128E",
X"1194",
X"128E",
X"130B",
X"1388",
X"1117",
X"1211",
X"1194",
X"1211",
X"109A",
X"0F23",
X"0DAC",
X"0CB2",
X"0947",
X"05DC",
X"02EE",
X"01F4",
X"0465",
X"02EE",
X"03E8",
X"0000",
X"0177",
X"FE89",
X"FB1E",
X"FB1E",
X"FE0C",
X"F9A7",
X"F8AD",
X"F830",
X"F448",
X"F63C",
X"F4C5",
X"F34E",
X"EF66",
X"EEE9",
X"F15A",
X"EE6C",
X"ED72",
X"EB01",
X"EA84",
X"EBFB",
X"ECF5",
X"ED72",
X"ECF5",
X"EEE9",
X"EF66",
X"F0DD",
X"F15A",
X"F2D1",
X"F3CB",
X"F448",
X"F15A",
X"F0DD",
X"F4C5",
X"F060",
X"F2D1",
X"F34E",
X"F3CB",
X"F7B3",
X"F542",
X"F92A",
X"FD12",
X"FB1E",
X"FC18",
X"FC18",
X"FA24",
X"FAA1",
X"F8AD",
X"F7B3",
X"F830",
X"F7B3",
X"F3CB",
X"F254",
X"ED72",
X"ED72",
X"F254",
X"F254",
X"F254",
X"EFE3",
X"F15A",
X"F15A",
X"EEE9",
X"EEE9",
X"EF66",
X"F060",
X"EE6C",
X"EEE9",
X"EE6C",
X"ED72",
X"ECF5",
X"EE6C",
X"EC78",
X"EB7E",
X"EC78",
X"E890",
X"EA07",
X"E61F",
X"E796",
X"EA84",
X"E98A",
X"EB01",
X"E890",
X"E813",
X"EBFB",
X"E98A",
X"E90D",
X"E98A",
X"EBFB",
X"ECF5",
X"ED72",
X"EEE9",
X"EFE3",
X"EEE9",
X"EEE9",
X"F0DD",
X"ED72",
X"F15A",
X"F2D1",
X"EFE3",
X"F254",
X"F1D7",
X"F2D1",
X"F3CB",
X"F1D7",
X"F060",
X"F3CB",
X"F542",
X"F542",
X"F736",
X"F6B9",
X"F830",
X"FAA1",
X"FC95",
X"0000",
X"00FA",
X"01F4",
X"02EE",
X"0465",
X"04E2",
X"0659",
X"0753",
X"04E2",
X"02EE",
X"02EE",
X"01F4",
X"01F4",
X"0177",
X"0271",
X"04E2",
X"04E2",
X"06D6",
X"06D6",
X"08CA",
X"0ABE",
X"0BB8",
X"0BB8",
X"0ABE",
X"0C35",
X"0C35",
X"0BB8",
X"0B3B",
X"0ABE",
X"0A41",
X"0A41",
X"08CA",
X"084D",
X"084D",
X"0947",
X"0ABE",
X"0947",
X"09C4",
X"0947",
X"0ABE",
X"0C35",
X"0B3B",
X"09C4",
X"08CA",
X"09C4",
X"0A41",
X"0947",
X"084D",
X"07D0",
X"06D6",
X"0947",
X"084D",
X"07D0",
X"09C4",
X"09C4",
X"0947",
X"09C4",
X"07D0",
X"09C4",
X"0947",
X"07D0",
X"0753",
X"08CA",
X"084D",
X"0753",
X"09C4",
X"0BB8",
X"0D2F",
X"0ABE",
X"0FA0",
X"0EA6",
X"0CB2",
X"101D",
X"0C35",
X"0EA6",
X"0D2F",
X"0CB2",
X"0D2F",
X"128E",
X"0E29",
X"0D2F",
X"1117",
X"0F23",
X"109A",
X"1117",
X"1482",
X"130B",
X"15F9",
X"15F9",
X"18E7",
X"16F3",
X"16F3",
X"1770",
X"15F9",
X"15F9",
X"1676",
X"1482",
X"15F9",
X"18E7",
X"186A",
X"16F3",
X"16F3",
X"1405",
X"16F3",
X"1211",
X"16F3",
X"1211",
X"1194",
X"130B",
X"0CB2",
X"0C35",
X"0C35",
X"0A41",
X"0B3B",
X"08CA",
X"07D0",
X"0659",
X"05DC",
X"04E2",
X"05DC",
X"03E8",
X"04E2",
X"0659",
X"0659",
X"0465",
X"06D6",
X"055F",
X"055F",
X"06D6",
X"055F",
X"04E2",
X"055F",
X"06D6",
X"04E2",
X"036B",
X"0465",
X"04E2",
X"036B",
X"036B",
X"0177",
X"0177",
X"FF83",
X"FF83",
X"00FA",
X"007D",
X"FD12",
X"FC95",
X"FD12",
X"FA24",
X"FAA1",
X"FB1E",
X"FB1E",
X"FC18",
X"FB9B",
X"F8AD",
X"F63C",
X"F7B3",
X"F8AD",
X"F830",
X"FA24",
X"F830",
X"F542",
X"F92A",
X"F34E",
X"F4C5",
X"F2D1",
X"F3CB",
X"F254",
X"F3CB",
X"F3CB",
X"F0DD",
X"F3CB",
X"F15A",
X"F448",
X"F448",
X"F2D1",
X"F3CB",
X"F1D7",
X"F15A",
X"F2D1",
X"F6B9",
X"F63C",
X"F6B9",
X"F542",
X"F6B9",
X"F63C",
X"F8AD",
X"F9A7",
X"F6B9",
X"F6B9",
X"F3CB",
X"F448",
X"F1D7",
X"F15A",
X"EEE9",
X"F15A",
X"F2D1",
X"EF66",
X"EF66",
X"ED72",
X"EEE9",
X"EF66",
X"EFE3",
X"F1D7",
X"F15A",
X"F0DD",
X"EEE9",
X"EDEF",
X"EE6C",
X"ECF5",
X"EA84",
X"E90D",
X"E719",
X"E69C",
X"E4A8",
X"E331",
X"E525",
X"E4A8",
X"E2B4",
X"E331",
X"E5A2",
X"E61F",
X"E42B",
X"E61F",
X"E719",
X"E4A8",
X"E5A2",
X"E69C",
X"E890",
X"EA07",
X"E890",
X"ECF5",
X"EB7E",
X"EC78",
X"F060",
X"F0DD",
X"EEE9",
X"F0DD",
X"F254",
X"F2D1",
X"F542",
X"F830",
X"F92A",
X"F8AD",
X"FB1E",
X"FD8F",
X"FE0C",
X"FE0C",
X"00FA",
X"0177",
X"0177",
X"01F4",
X"02EE",
X"0177",
X"01F4",
X"0659",
X"0753",
X"07D0",
X"084D",
X"084D",
X"0947",
X"0ABE",
X"0B3B",
X"0ABE",
X"09C4",
X"0947",
X"07D0",
X"05DC",
X"05DC",
X"055F",
X"055F",
X"055F",
X"0659",
X"06D6",
X"0753",
X"06D6",
X"0659",
X"0659",
X"0465",
X"02EE",
X"00FA",
X"007D",
X"FF83",
X"FE89",
X"FE89",
X"FE0C",
X"FD12",
X"FC95",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE89",
X"0000",
X"FF83",
X"00FA",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"02EE",
X"04E2",
X"03E8",
X"04E2",
X"05DC",
X"06D6",
X"06D6",
X"06D6",
X"0947",
X"0B3B",
X"0BB8",
X"0B3B",
X"0BB8",
X"0D2F",
X"0DAC",
X"0EA6",
X"0FA0",
X"1211",
X"128E",
X"1405",
X"16F3",
X"1770",
X"1770",
X"1676",
X"1770",
X"17ED",
X"186A",
X"19E1",
X"1964",
X"19E1",
X"1B58",
X"1CCF",
X"1C52",
X"1E46",
X"1C52",
X"1C52",
X"1DC9",
X"1E46",
X"20B7",
X"1FBD",
X"1F40",
X"1CCF",
X"1CCF",
X"1BD5",
X"1ADB",
X"18E7",
X"18E7",
X"1BD5",
X"1E46",
X"1CCF",
X"1A5E",
X"18E7",
X"18E7",
X"19E1",
X"1A5E",
X"1ADB",
X"18E7",
X"14FF",
X"128E",
X"1405",
X"157C",
X"1194",
X"0F23",
X"101D",
X"0F23",
X"0B3B",
X"07D0",
X"03E8",
X"02EE",
X"03E8",
X"01F4",
X"00FA",
X"01F4",
X"0177",
X"FE0C",
X"FAA1",
X"FB9B",
X"FB1E",
X"F8AD",
X"F5BF",
X"F736",
X"F7B3",
X"F736",
X"F63C",
X"F5BF",
X"F542",
X"F4C5",
X"F5BF",
X"F63C",
X"F4C5",
X"F448",
X"F7B3",
X"F6B9",
X"F34E",
X"F34E",
X"F448",
X"F4C5",
X"F254",
X"F15A",
X"F15A",
X"F2D1",
X"F34E",
X"F1D7",
X"F34E",
X"F5BF",
X"F5BF",
X"F736",
X"F736",
X"F830",
X"F4C5",
X"F1D7",
X"F34E",
X"F15A",
X"F15A",
X"EE6C",
X"F0DD",
X"EF66",
X"EC78",
X"ECF5",
X"EE6C",
X"EE6C",
X"EF66",
X"ECF5",
X"EB7E",
X"EDEF",
X"EE6C",
X"EE6C",
X"EBFB",
X"EBFB",
X"EC78",
X"E98A",
X"E890",
X"EB01",
X"EA07",
X"E796",
X"E890",
X"EBFB",
X"ED72",
X"EEE9",
X"EFE3",
X"EF66",
X"EEE9",
X"EEE9",
X"F0DD",
X"F1D7",
X"F0DD",
X"F15A",
X"F2D1",
X"F254",
X"F2D1",
X"F3CB",
X"F254",
X"F2D1",
X"F542",
X"F92A",
X"FAA1",
X"FA24",
X"FB1E",
X"FB9B",
X"FA24",
X"FC95",
X"FE0C",
X"FF83",
X"03E8",
X"01F4",
X"0271",
X"0271",
X"0465",
X"0753",
X"04E2",
X"03E8",
X"02EE",
X"04E2",
X"055F",
X"055F",
X"06D6",
X"07D0",
X"084D",
X"08CA",
X"09C4",
X"084D",
X"084D",
X"08CA",
X"0753",
X"0465",
X"0465",
X"0465",
X"02EE",
X"007D",
X"007D",
X"00FA",
X"0271",
X"0659",
X"07D0",
X"036B",
X"0271",
X"0465",
X"0659",
X"03E8",
X"03E8",
X"04E2",
X"01F4",
X"0177",
X"01F4",
X"036B",
X"01F4",
X"0271",
X"0271",
X"0271",
X"036B",
X"0465",
X"03E8",
X"03E8",
X"036B",
X"04E2",
X"055F",
X"04E2",
X"036B",
X"0000",
X"0465",
X"05DC",
X"03E8",
X"007D",
X"01F4",
X"0271",
X"0000",
X"FF06",
X"FE89",
X"FE89",
X"FD12",
X"FD8F",
X"FC18",
X"FC18",
X"FD12",
X"FB1E",
X"F8AD",
X"F8AD",
X"F8AD",
X"F736",
X"F7B3",
X"F8AD",
X"F8AD",
X"F736",
X"F7B3",
X"F6B9",
X"F5BF",
X"F736",
X"F5BF",
X"F448",
X"F2D1",
X"F448",
X"F4C5",
X"F63C",
X"F7B3",
X"F92A",
X"FAA1",
X"FD12",
X"FF83",
X"007D",
X"00FA",
X"00FA",
X"01F4",
X"02EE",
X"036B",
X"03E8",
X"0465",
X"03E8",
X"03E8",
X"03E8",
X"02EE",
X"02EE",
X"03E8",
X"03E8",
X"0465",
X"036B",
X"0271",
X"0271",
X"055F",
X"06D6",
X"0753",
X"08CA",
X"0A41",
X"0CB2",
X"0A41",
X"08CA",
X"09C4",
X"08CA",
X"084D",
X"07D0",
X"084D",
X"0753",
X"07D0",
X"08CA",
X"0659",
X"0465",
X"04E2",
X"07D0",
X"0659",
X"05DC",
X"07D0",
X"0947",
X"09C4",
X"06D6",
X"04E2",
X"02EE",
X"0000",
X"0000",
X"01F4",
X"00FA",
X"01F4",
X"00FA",
X"007D",
X"0000",
X"007D",
X"FE0C",
X"FE0C",
X"0271",
X"01F4",
X"03E8",
X"036B",
X"01F4",
X"036B",
X"03E8",
X"03E8",
X"036B",
X"036B",
X"07D0",
X"04E2",
X"055F",
X"03E8",
X"06D6",
X"04E2",
X"0753",
X"04E2",
X"0ABE",
X"05DC",
X"0947",
X"08CA",
X"0A41",
X"0B3B",
X"0C35",
X"0947",
X"09C4",
X"09C4",
X"09C4",
X"0DAC",
X"0A41",
X"0ABE",
X"0947",
X"055F",
X"06D6",
X"055F",
X"084D",
X"0753",
X"084D",
X"07D0",
X"0BB8",
X"0753",
X"09C4",
X"0753",
X"0465",
X"05DC",
X"036B",
X"0177",
X"0271",
X"01F4",
X"007D",
X"0271",
X"007D",
X"0000",
X"007D",
X"0000",
X"02EE",
X"FD8F",
X"0000",
X"036B",
X"01F4",
X"0271",
X"036B",
X"0271",
X"036B",
X"02EE",
X"0465",
X"007D",
X"007D",
X"0271",
X"01F4",
X"FE89",
X"FD8F",
X"FD8F",
X"FD12",
X"FC95",
X"FB1E",
X"FB9B",
X"FB9B",
X"FA24",
X"F7B3",
X"F34E",
X"F3CB",
X"F8AD",
X"F8AD",
X"F830",
X"F63C",
X"F63C",
X"F542",
X"F2D1",
X"F254",
X"F2D1",
X"F15A",
X"F3CB",
X"F6B9",
X"FB1E",
X"F8AD",
X"F6B9",
X"F9A7",
X"FA24",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FF06",
X"00FA",
X"02EE",
X"007D",
X"007D",
X"036B",
X"007D",
X"FE89",
X"FF83",
X"FC95",
X"FF83",
X"03E8",
X"05DC",
X"06D6",
X"05DC",
X"06D6",
X"06D6",
X"0753",
X"055F",
X"0177",
X"0000",
X"FE0C",
X"FC18",
X"FE0C",
X"007D",
X"00FA",
X"0000",
X"FF83",
X"FF06",
X"FB9B",
X"F830",
X"F6B9",
X"F7B3",
X"FD12",
X"FF06",
X"FE0C",
X"FC95",
X"FA24",
X"F92A",
X"F5BF",
X"F4C5",
X"F736",
X"F736",
X"F6B9",
X"F6B9",
X"F5BF",
X"F542",
X"F63C",
X"F736",
X"F5BF",
X"F6B9",
X"F63C",
X"F63C",
X"F34E",
X"F5BF",
X"F8AD",
X"F6B9",
X"F830",
X"F830",
X"F8AD",
X"F92A",
X"F7B3",
X"FB1E",
X"F92A",
X"F830",
X"F830",
X"F6B9",
X"F7B3",
X"F7B3",
X"F830",
X"F830",
X"F7B3",
X"F8AD",
X"F92A",
X"F5BF",
X"F5BF",
X"F5BF",
X"F6B9",
X"F7B3",
X"FA24",
X"FAA1",
X"FA24",
X"F8AD",
X"F92A",
X"FAA1",
X"FB1E",
X"FB1E",
X"FC95",
X"FE0C",
X"FE89",
X"FE89",
X"FD12",
X"FE0C",
X"FF83",
X"007D",
X"0271",
X"007D",
X"007D",
X"00FA",
X"0177",
X"02EE",
X"0177",
X"0177",
X"00FA",
X"FF06",
X"FE0C",
X"FF83",
X"007D",
X"0177",
X"02EE",
X"007D",
X"007D",
X"0177",
X"007D",
X"FF83",
X"00FA",
X"0271",
X"03E8",
X"0465",
X"055F",
X"055F",
X"0659",
X"06D6",
X"055F",
X"0465",
X"036B",
X"0271",
X"02EE",
X"02EE",
X"036B",
X"0271",
X"01F4",
X"007D",
X"0271",
X"036B",
X"036B",
X"01F4",
X"036B",
X"0177",
X"FE0C",
X"FF06",
X"FF06",
X"0177",
X"FE89",
X"FC95",
X"FF83",
X"FD12",
X"FC95",
X"FD12",
X"FF06",
X"007D",
X"0000",
X"0000",
X"00FA",
X"0177",
X"0000",
X"0271",
X"0177",
X"00FA",
X"01F4",
X"01F4",
X"02EE",
X"03E8",
X"02EE",
X"036B",
X"04E2",
X"04E2",
X"06D6",
X"055F",
X"0465",
X"04E2",
X"0659",
X"05DC",
X"055F",
X"05DC",
X"0753",
X"06D6",
X"05DC",
X"036B",
X"0465",
X"04E2",
X"05DC",
X"06D6",
X"07D0",
X"084D",
X"09C4",
X"0947",
X"0B3B",
X"0A41",
X"09C4",
X"0DAC",
X"0947",
X"0ABE",
X"0BB8",
X"0ABE",
X"0ABE",
X"0A41",
X"0BB8",
X"0A41",
X"0A41",
X"0BB8",
X"0C35",
X"0ABE",
X"0947",
X"0BB8",
X"0BB8",
X"0A41",
X"09C4",
X"0ABE",
X"0A41",
X"0A41",
X"0ABE",
X"0B3B",
X"0CB2",
X"0C35",
X"0D2F",
X"0CB2",
X"0DAC",
X"0EA6",
X"0E29",
X"0EA6",
X"0DAC",
X"0C35",
X"0C35",
X"0CB2",
X"0CB2",
X"0D2F",
X"0CB2",
X"0B3B",
X"0A41",
X"084D",
X"07D0",
X"0753",
X"084D",
X"0947",
X"09C4",
X"0A41",
X"0A41",
X"09C4",
X"08CA",
X"0753",
X"0659",
X"0659",
X"06D6",
X"0753",
X"0465",
X"036B",
X"0659",
X"0659",
X"0271",
X"02EE",
X"02EE",
X"036B",
X"055F",
X"03E8",
X"0177",
X"00FA",
X"007D",
X"FF06",
X"FD12",
X"FC95",
X"FC18",
X"FAA1",
X"F6B9",
X"F5BF",
X"F4C5",
X"F2D1",
X"F1D7",
X"EFE3",
X"EF66",
X"F060",
X"EE6C",
X"EE6C",
X"EE6C",
X"EBFB",
X"EB01",
X"EA84",
X"EB7E",
X"EBFB",
X"EB7E",
X"EB01",
X"EBFB",
X"EA84",
X"EBFB",
X"ECF5",
X"EDEF",
X"EFE3",
X"F1D7",
X"F254",
X"F254",
X"F3CB",
X"F542",
X"F5BF",
X"F6B9",
X"F830",
X"F8AD",
X"FAA1",
X"FA24",
X"FB1E",
X"FB9B",
X"FD12",
X"FB1E",
X"FC95",
X"FE0C",
X"FD12",
X"FC95",
X"FC18",
X"FB9B",
X"FA24",
X"FB1E",
X"F92A",
X"FA24",
X"F9A7",
X"F9A7",
X"F92A",
X"F830",
X"F830",
X"F7B3",
X"F8AD",
X"F830",
X"F8AD",
X"F736",
X"F63C",
X"F63C",
X"F542",
X"F34E",
X"F1D7",
X"F254",
X"F15A",
X"F1D7",
X"F34E",
X"F1D7",
X"F254",
X"F1D7",
X"F254",
X"F0DD",
X"F2D1",
X"F3CB",
X"F1D7",
X"F4C5",
X"F5BF",
X"F5BF",
X"F4C5",
X"F4C5",
X"F448",
X"F542",
X"F5BF",
X"F5BF",
X"F736",
X"F63C",
X"F92A",
X"F9A7",
X"F92A",
X"FB1E",
X"FB9B",
X"FB9B",
X"FD12",
X"FF06",
X"FF06",
X"007D",
X"0177",
X"00FA",
X"01F4",
X"03E8",
X"03E8",
X"04E2",
X"05DC",
X"0659",
X"05DC",
X"036B",
X"06D6",
X"055F",
X"05DC",
X"06D6",
X"05DC",
X"0659",
X"05DC",
X"06D6",
X"05DC",
X"05DC",
X"04E2",
X"0659",
X"0659",
X"04E2",
X"05DC",
X"05DC",
X"03E8",
X"0465",
X"055F",
X"04E2",
X"0659",
X"07D0",
X"07D0",
X"08CA",
X"08CA",
X"084D",
X"07D0",
X"06D6",
X"0659",
X"06D6",
X"05DC",
X"055F",
X"055F",
X"0465",
X"0465",
X"036B",
X"0271",
X"01F4",
X"0271",
X"0177",
X"02EE",
X"036B",
X"00FA",
X"036B",
X"036B",
X"0271",
X"036B",
X"0465",
X"0465",
X"0465",
X"0659",
X"05DC",
X"0753",
X"0659",
X"05DC",
X"07D0",
X"084D",
X"06D6",
X"05DC",
X"07D0",
X"07D0",
X"0753",
X"0753",
X"07D0",
X"0753",
X"07D0",
X"07D0",
X"08CA",
X"0947",
X"06D6",
X"07D0",
X"084D",
X"0659",
X"084D",
X"0947",
X"0947",
X"0947",
X"08CA",
X"07D0",
X"0753",
X"0659",
X"0465",
X"0465",
X"055F",
X"04E2",
X"03E8",
X"03E8",
X"0465",
X"036B",
X"0465",
X"04E2",
X"03E8",
X"02EE",
X"0271",
X"01F4",
X"0177",
X"00FA",
X"00FA",
X"0177",
X"00FA",
X"0177",
X"00FA",
X"007D",
X"0177",
X"0177",
X"0177",
X"0271",
X"036B",
X"036B",
X"04E2",
X"05DC",
X"04E2",
X"05DC",
X"0659",
X"0659",
X"06D6",
X"05DC",
X"0659",
X"0753",
X"06D6",
X"0753",
X"0753",
X"07D0",
X"08CA",
X"08CA",
X"09C4",
X"09C4",
X"0ABE",
X"0A41",
X"0B3B",
X"0ABE",
X"0B3B",
X"09C4",
X"08CA",
X"08CA",
X"084D",
X"0659",
X"05DC",
X"05DC",
X"04E2",
X"04E2",
X"0465",
X"03E8",
X"036B",
X"02EE",
X"036B",
X"03E8",
X"0465",
X"036B",
X"02EE",
X"036B",
X"0271",
X"00FA",
X"FF83",
X"FF06",
X"FE89",
X"FE89",
X"FE0C",
X"FD12",
X"FD12",
X"FD12",
X"FC18",
X"FC95",
X"FC95",
X"FC95",
X"FD12",
X"FD8F",
X"FE0C",
X"FE89",
X"FD8F",
X"FE0C",
X"FF06",
X"FF83",
X"0000",
X"FE0C",
X"FF06",
X"FF06",
X"FF06",
X"FE89",
X"FD8F",
X"FD8F",
X"FE89",
X"FD8F",
X"FD8F",
X"FE89",
X"FC95",
X"FD8F",
X"FC18",
X"FAA1",
X"FC18",
X"FB1E",
X"F8AD",
X"F736",
X"F736",
X"F736",
X"F5BF",
X"F542",
X"F448",
X"F34E",
X"F254",
X"F1D7",
X"F15A",
X"F060",
X"F060",
X"F060",
X"EFE3",
X"EEE9",
X"EE6C",
X"EE6C",
X"EDEF",
X"ED72",
X"ED72",
X"ED72",
X"EDEF",
X"EDEF",
X"EEE9",
X"EEE9",
X"EE6C",
X"EEE9",
X"EE6C",
X"EDEF",
X"ED72",
X"EC78",
X"EC78",
X"EC78",
X"EE6C",
X"EF66",
X"EEE9",
X"EEE9",
X"F060",
X"EFE3",
X"F0DD",
X"F15A",
X"F15A",
X"F2D1",
X"F254",
X"F0DD",
X"F0DD",
X"F15A",
X"F254",
X"F2D1",
X"F254",
X"F34E",
X"F3CB",
X"F3CB",
X"F448",
X"F6B9",
X"F63C",
X"F63C",
X"F7B3",
X"F736",
X"F736",
X"F830",
X"F830",
X"F7B3",
X"FA24",
X"FA24",
X"FA24",
X"FAA1",
X"FD12",
X"FD8F",
X"FD8F",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"00FA",
X"007D",
X"007D",
X"0271",
X"036B",
X"03E8",
X"0465",
X"04E2",
X"0659",
X"05DC",
X"0659",
X"0659",
X"0659",
X"0753",
X"08CA",
X"0947",
X"09C4",
X"0A41",
X"0947",
X"09C4",
X"0ABE",
X"0C35",
X"0CB2",
X"0B3B",
X"09C4",
X"0B3B",
X"0BB8",
X"0BB8",
X"0C35",
X"0CB2",
X"0D2F",
X"0DAC",
X"0D2F",
X"0D2F",
X"0D2F",
X"0F23",
X"0F23",
X"0FA0",
X"101D",
X"101D",
X"109A",
X"109A",
X"109A",
X"0FA0",
X"0FA0",
X"0EA6",
X"0F23",
X"101D",
X"109A",
X"1117",
X"1117",
X"1194",
X"1211",
X"130B",
X"130B",
X"1482",
X"1482",
X"1388",
X"1388",
X"130B",
X"1211",
X"1117",
X"1117",
X"101D",
X"101D",
X"101D",
X"101D",
X"0FA0",
X"0F23",
X"0E29",
X"0DAC",
X"0E29",
X"0E29",
X"0DAC",
X"0D2F",
X"0CB2",
X"0BB8",
X"0BB8",
X"0C35",
X"09C4",
X"07D0",
X"0753",
X"0753",
X"055F",
X"055F",
X"0465",
X"036B",
X"0465",
X"03E8",
X"0465",
X"036B",
X"0271",
X"01F4",
X"007D",
X"00FA",
X"FF83",
X"FE89",
X"0000",
X"FF06",
X"FE0C",
X"FD12",
X"FE89",
X"FD8F",
X"FC95",
X"FB9B",
X"FAA1",
X"FB1E",
X"FC18",
X"FC95",
X"FD8F",
X"FE89",
X"FE89",
X"FE0C",
X"FD8F",
X"FE0C",
X"FE0C",
X"FD12",
X"FD8F",
X"FE89",
X"FF06",
X"FD12",
X"FD12",
X"FD8F",
X"FC95",
X"FC95",
X"FD12",
X"FC95",
X"FC18",
X"FD12",
X"FD8F",
X"FC18",
X"FB9B",
X"FB1E",
X"FC18",
X"FB9B",
X"FA24",
X"FA24",
X"F9A7",
X"F830",
X"F6B9",
X"F736",
X"F830",
X"F92A",
X"F736",
X"F7B3",
X"F7B3",
X"F8AD",
X"F8AD",
X"F6B9",
X"F7B3",
X"F736",
X"F736",
X"F7B3",
X"F736",
X"F63C",
X"F736",
X"F7B3",
X"F830",
X"F830",
X"F736",
X"F830",
X"F92A",
X"F9A7",
X"F9A7",
X"F9A7",
X"FB1E",
X"FA24",
X"F9A7",
X"FAA1",
X"F8AD",
X"F8AD",
X"F830",
X"F6B9",
X"F6B9",
X"F542",
X"F542",
X"F542",
X"F448",
X"F448",
X"F63C",
X"F63C",
X"F63C",
X"F5BF",
X"F6B9",
X"F542",
X"F3CB",
X"F448",
X"F254",
X"F34E",
X"F254",
X"F15A",
X"F1D7",
X"F15A",
X"EEE9",
X"EEE9",
X"EE6C",
X"EE6C",
X"F060",
X"EFE3",
X"F15A",
X"F2D1",
X"F1D7",
X"F448",
X"F4C5",
X"F4C5",
X"F5BF",
X"F63C",
X"F6B9",
X"F5BF",
X"F92A",
X"FAA1",
X"FB9B",
X"FC95",
X"FE89",
X"0000",
X"0000",
X"007D",
X"00FA",
X"01F4",
X"036B",
X"055F",
X"05DC",
X"084D",
X"07D0",
X"07D0",
X"07D0",
X"08CA",
X"0753",
X"08CA",
X"08CA",
X"08CA",
X"0947",
X"084D",
X"084D",
X"08CA",
X"09C4",
X"084D",
X"08CA",
X"0947",
X"07D0",
X"07D0",
X"084D",
X"07D0",
X"07D0",
X"07D0",
X"06D6",
X"084D",
X"07D0",
X"0753",
X"05DC",
X"05DC",
X"055F",
X"03E8",
X"04E2",
X"03E8",
X"055F",
X"036B",
X"0271",
X"01F4",
X"01F4",
X"0000",
X"FE89",
X"FE0C",
X"FD8F",
X"FE0C",
X"FF06",
X"0000",
X"FE0C",
X"FF83",
X"0000",
X"FE0C",
X"FF06",
X"FE0C",
X"FE0C",
X"FE89",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE89",
X"FF06",
X"FE89",
X"0000",
X"01F4",
X"0177",
X"0000",
X"02EE",
X"036B",
X"0465",
X"04E2",
X"055F",
X"05DC",
X"0659",
X"0465",
X"04E2",
X"055F",
X"055F",
X"0753",
X"0753",
X"07D0",
X"084D",
X"084D",
X"084D",
X"0A41",
X"0BB8",
X"0ABE",
X"0B3B",
X"0C35",
X"0ABE",
X"0A41",
X"0947",
X"09C4",
X"08CA",
X"084D",
X"0947",
X"08CA",
X"0753",
X"0753",
X"07D0",
X"0753",
X"0753",
X"05DC",
X"055F",
X"0465",
X"036B",
X"0271",
X"01F4",
X"0271",
X"01F4",
X"01F4",
X"00FA",
X"FF06",
X"FE89",
X"FF06",
X"FF83",
X"FE0C",
X"FD12",
X"FD8F",
X"FD12",
X"FB1E",
X"FB9B",
X"FB1E",
X"FAA1",
X"FAA1",
X"FB9B",
X"FB1E",
X"FB9B",
X"FD8F",
X"FD8F",
X"FE0C",
X"FD12",
X"FE0C",
X"FF06",
X"FF06",
X"FF06",
X"FE0C",
X"FF06",
X"FE89",
X"FF06",
X"0000",
X"0000",
X"007D",
X"00FA",
X"FF83",
X"007D",
X"01F4",
X"0271",
X"02EE",
X"01F4",
X"036B",
X"0271",
X"0271",
X"0271",
X"01F4",
X"02EE",
X"02EE",
X"04E2",
X"04E2",
X"04E2",
X"05DC",
X"05DC",
X"055F",
X"0659",
X"06D6",
X"04E2",
X"0465",
X"055F",
X"036B",
X"02EE",
X"0271",
X"01F4",
X"02EE",
X"036B",
X"03E8",
X"01F4",
X"036B",
X"036B",
X"0271",
X"03E8",
X"01F4",
X"0177",
X"02EE",
X"01F4",
X"0271",
X"00FA",
X"007D",
X"0000",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE0C",
X"FD12",
X"FD12",
X"FB1E",
X"FB1E",
X"FB9B",
X"FA24",
X"FB1E",
X"F8AD",
X"F736",
X"F63C",
X"F5BF",
X"F542",
X"F4C5",
X"F5BF",
X"F6B9",
X"F6B9",
X"F4C5",
X"F542",
X"F63C",
X"F63C",
X"F542",
X"F542",
X"F5BF",
X"F542",
X"F2D1",
X"F542",
X"F542",
X"F4C5",
X"F63C",
X"F830",
X"F6B9",
X"F542",
X"F736",
X"F6B9",
X"F7B3",
X"F736",
X"F6B9",
X"F7B3",
X"F92A",
X"F830",
X"F8AD",
X"F9A7",
X"F830",
X"F830",
X"FB9B",
X"FA24",
X"FA24",
X"FC18",
X"FB1E",
X"FC95",
X"FC95",
X"FB9B",
X"FC18",
X"FC18",
X"FE89",
X"FF83",
X"FB9B",
X"FF06",
X"0000",
X"FD12",
X"FE89",
X"FF06",
X"FD12",
X"FE0C",
X"FE0C",
X"FB1E",
X"FC95",
X"FE0C",
X"FF06",
X"0000",
X"007D",
X"02EE",
X"02EE",
X"01F4",
X"01F4",
X"0177",
X"00FA",
X"00FA",
X"01F4",
X"0271",
X"01F4",
X"0271",
X"02EE",
X"02EE",
X"03E8",
X"03E8",
X"0271",
X"03E8",
X"03E8",
X"01F4",
X"0271",
X"03E8",
X"04E2",
X"055F",
X"05DC",
X"055F",
X"03E8",
X"0465",
X"05DC",
X"0465",
X"04E2",
X"0753",
X"06D6",
X"0659",
X"04E2",
X"04E2",
X"0753",
X"07D0",
X"055F",
X"05DC",
X"0659",
X"0753",
X"06D6",
X"0753",
X"0753",
X"07D0",
X"06D6",
X"0659",
X"06D6",
X"0753",
X"06D6",
X"06D6",
X"084D",
X"0947",
X"084D",
X"07D0",
X"0947",
X"07D0",
X"084D",
X"08CA",
X"084D",
X"0947",
X"09C4",
X"0753",
X"06D6",
X"07D0",
X"0947",
X"07D0",
X"0659",
X"05DC",
X"0465",
X"055F",
X"06D6",
X"055F",
X"04E2",
X"05DC",
X"0659",
X"04E2",
X"055F",
X"055F",
X"055F",
X"0465",
X"03E8",
X"0271",
X"01F4",
X"0177",
X"FF06",
X"FE0C",
X"FE0C",
X"FD12",
X"FC95",
X"FB9B",
X"FB9B",
X"FB1E",
X"FAA1",
X"FB9B",
X"FB9B",
X"FC18",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC95",
X"FC95",
X"FD12",
X"FD8F",
X"FE0C",
X"FE0C",
X"FD12",
X"FD12",
X"FD12",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FE0C",
X"FD12",
X"FD12",
X"FD8F",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FD12",
X"FC95",
X"FC95",
X"FC18",
X"FC95",
X"FC95",
X"FB9B",
X"FC95",
X"FD12",
X"FC18",
X"FC18",
X"FD12",
X"FD12",
X"FC95",
X"FE0C",
X"FE0C",
X"FD12",
X"FE0C",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"FE89",
X"FE0C",
X"FE89",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FD8F",
X"FD8F",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"FF83",
X"0000",
X"FF06",
X"FD8F",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD12",
X"FE89",
X"FF83",
X"FF06",
X"FE0C",
X"FD8F",
X"FD12",
X"FE0C",
X"FE89",
X"FE89",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD12",
X"FC95",
X"FC18",
X"FB9B",
X"FB9B",
X"FC18",
X"FB9B",
X"FB1E",
X"FB9B",
X"FB9B",
X"FC18",
X"FC18",
X"FC18",
X"FB9B",
X"FC18",
X"FD12",
X"FC95",
X"FD12",
X"FD8F",
X"FC95",
X"FC18",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FE89",
X"FF06",
X"FD12",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE0C",
X"FD8F",
X"FE0C",
X"FD8F",
X"FD12",
X"FB1E",
X"FB9B",
X"FD12",
X"FC18",
X"FAA1",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB1E",
X"FAA1",
X"FB9B",
X"FB1E",
X"FB9B",
X"FB9B",
X"FAA1",
X"FB1E",
X"FD8F",
X"FE89",
X"FD8F",
X"FE89",
X"FE0C",
X"FF83",
X"00FA",
X"FF06",
X"007D",
X"01F4",
X"00FA",
X"01F4",
X"0465",
X"04E2",
X"04E2",
X"0465",
X"055F",
X"05DC",
X"0753",
X"06D6",
X"05DC",
X"07D0",
X"0659",
X"04E2",
X"05DC",
X"07D0",
X"08CA",
X"0753",
X"055F",
X"0753",
X"07D0",
X"0659",
X"0659",
X"06D6",
X"0659",
X"05DC",
X"04E2",
X"055F",
X"05DC",
X"055F",
X"0753",
X"06D6",
X"0753",
X"084D",
X"05DC",
X"06D6",
X"0659",
X"06D6",
X"06D6",
X"0659",
X"05DC",
X"0753",
X"07D0",
X"07D0",
X"07D0",
X"0947",
X"0ABE",
X"0A41",
X"09C4",
X"09C4",
X"09C4",
X"0A41",
X"09C4",
X"0947",
X"0947",
X"08CA",
X"084D",
X"084D",
X"07D0",
X"0659",
X"0659",
X"0659",
X"08CA",
X"09C4",
X"084D",
X"0659",
X"0659",
X"05DC",
X"05DC",
X"04E2",
X"04E2",
X"03E8",
X"0271",
X"0465",
X"055F",
X"0271",
X"00FA",
X"036B",
X"01F4",
X"0000",
X"00FA",
X"03E8",
X"02EE",
X"FF83",
X"01F4",
X"01F4",
X"0000",
X"00FA",
X"00FA",
X"00FA",
X"0177",
X"007D",
X"FF06",
X"FF83",
X"007D",
X"007D",
X"0000",
X"FE89",
X"FD8F",
X"FF06",
X"0000",
X"FE0C",
X"FB1E",
X"FB9B",
X"FD12",
X"FE89",
X"FC95",
X"FB9B",
X"FD12",
X"FB1E",
X"FAA1",
X"FB1E",
X"FAA1",
X"FA24",
X"F9A7",
X"FA24",
X"F9A7",
X"F7B3",
X"F7B3",
X"F7B3",
X"F63C",
X"F830",
X"F8AD",
X"F5BF",
X"F448",
X"F5BF",
X"F5BF",
X"F542",
X"F5BF",
X"F5BF",
X"F736",
X"F63C",
X"F4C5",
X"F5BF",
X"F4C5",
X"F4C5",
X"F63C",
X"F736",
X"F5BF",
X"F736",
X"F830",
X"F6B9",
X"F63C",
X"F6B9",
X"F736",
X"F7B3",
X"F92A",
X"F8AD",
X"F8AD",
X"F92A",
X"F92A",
X"F9A7",
X"FA24",
X"F9A7",
X"F9A7",
X"FB9B",
X"FB9B",
X"FB1E",
X"FAA1",
X"FB9B",
X"FD8F",
X"FD8F",
X"FC18",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FD12",
X"FD8F",
X"FD8F",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"FF83",
X"0000",
X"007D",
X"FF83",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"01F4",
X"0177",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"00FA",
X"0177",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"0177",
X"00FA",
X"0177",
X"0271",
X"0177",
X"0177",
X"0271",
X"036B",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"00FA",
X"0177",
X"0177",
X"00FA",
X"FF83",
X"007D",
X"0000",
X"007D",
X"00FA",
X"007D",
X"0177",
X"00FA",
X"0177",
X"01F4",
X"0177",
X"0177",
X"0177",
X"01F4",
X"0177",
X"0177",
X"0177",
X"01F4",
X"0271",
X"0271",
X"036B",
X"03E8",
X"03E8",
X"0465",
X"04E2",
X"055F",
X"055F",
X"05DC",
X"05DC",
X"0659",
X"0659",
X"06D6",
X"0753",
X"0753",
X"07D0",
X"07D0",
X"07D0",
X"08CA",
X"0947",
X"0A41",
X"0A41",
X"0B3B",
X"0BB8",
X"0BB8",
X"0B3B",
X"0C35",
X"0C35",
X"0C35",
X"0BB8",
X"0B3B",
X"0B3B",
X"0B3B",
X"0B3B",
X"0ABE",
X"0ABE",
X"0B3B",
X"0ABE",
X"0ABE",
X"0B3B",
X"0A41",
X"0947",
X"09C4",
X"0947",
X"08CA",
X"084D",
X"07D0",
X"06D6",
X"055F",
X"04E2",
X"0465",
X"036B",
X"02EE",
X"01F4",
X"0177",
X"007D",
X"FF06",
X"FE89",
X"FD8F",
X"FD12",
X"FD8F",
X"FC18",
X"FB1E",
X"FAA1",
X"F9A7",
X"F8AD",
X"F8AD",
X"F8AD",
X"F830",
X"F736",
X"F6B9",
X"F736",
X"F6B9",
X"F63C",
X"F5BF",
X"F542",
X"F5BF",
X"F4C5",
X"F448",
X"F448",
X"F3CB",
X"F3CB",
X"F2D1",
X"F2D1",
X"F2D1",
X"F1D7",
X"F254",
X"F2D1",
X"F3CB",
X"F34E",
X"F1D7",
X"F254",
X"F34E",
X"F3CB",
X"F34E",
X"F3CB",
X"F542",
X"F5BF",
X"F6B9",
X"F736",
X"F736",
X"F830",
X"FA24",
X"FB1E",
X"FC18",
X"FC18",
X"FD12",
X"FE0C",
X"FE89",
X"FE0C",
X"FF83",
X"007D",
X"0000",
X"0000",
X"0000",
X"FF83",
X"00FA",
X"0000",
X"0000",
X"007D",
X"0000",
X"FF06",
X"0000",
X"007D",
X"0000",
X"007D",
X"007D",
X"0000",
X"FF06",
X"FF06",
X"FF83",
X"FE89",
X"FD8F",
X"FE89",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD12",
X"FC95",
X"FC95",
X"FD12",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0177",
X"00FA",
X"00FA",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"02EE",
X"03E8",
X"03E8",
X"04E2",
X"05DC",
X"05DC",
X"05DC",
X"0659",
X"07D0",
X"0753",
X"06D6",
X"0659",
X"06D6",
X"06D6",
X"0659",
X"0659",
X"0659",
X"055F",
X"05DC",
X"06D6",
X"06D6",
X"0659",
X"06D6",
X"0659",
X"0659",
X"0659",
X"04E2",
X"055F",
X"055F",
X"05DC",
X"05DC",
X"05DC",
X"055F",
X"05DC",
X"0659",
X"0659",
X"0659",
X"055F",
X"055F",
X"05DC",
X"05DC",
X"055F",
X"04E2",
X"055F",
X"04E2",
X"0465",
X"04E2",
X"055F",
X"0465",
X"055F",
X"055F",
X"055F",
X"0659",
X"055F",
X"055F",
X"05DC",
X"05DC",
X"04E2",
X"0465",
X"03E8",
X"03E8",
X"036B",
X"02EE",
X"01F4",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"036B",
X"0271",
X"0271",
X"0177",
X"0177",
X"01F4",
X"0177",
X"0271",
X"0177",
X"007D",
X"00FA",
X"0177",
X"007D",
X"0000",
X"007D",
X"007D",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FE0C",
X"FD8F",
X"FE0C",
X"FD8F",
X"FC95",
X"FD12",
X"FD12",
X"FC95",
X"FC18",
X"FB1E",
X"FB9B",
X"FB1E",
X"FA24",
X"FA24",
X"FA24",
X"FA24",
X"F8AD",
X"F9A7",
X"F92A",
X"F8AD",
X"F830",
X"F7B3",
X"F8AD",
X"F830",
X"F7B3",
X"F8AD",
X"F8AD",
X"F7B3",
X"F8AD",
X"F8AD",
X"F8AD",
X"F8AD",
X"F830",
X"F8AD",
X"F8AD",
X"F7B3",
X"F7B3",
X"F7B3",
X"F8AD",
X"F9A7",
X"F9A7",
X"F9A7",
X"FA24",
X"F9A7",
X"FAA1",
X"FB1E",
X"FB1E",
X"FB9B",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FD12",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"FF06",
X"FF06",
X"FF83",
X"FE89",
X"FF83",
X"0000",
X"007D",
X"007D",
X"0000",
X"007D",
X"0000",
X"007D",
X"0000",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF06",
X"FE89",
X"FE89",
X"FE0C",
X"FD8F",
X"FE0C",
X"FC95",
X"FC18",
X"FC18",
X"FC95",
X"FD12",
X"FC95",
X"FD12",
X"FD8F",
X"FC95",
X"FC18",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FC95",
X"FD12",
X"FD12",
X"FD8F",
X"FC95",
X"FD12",
X"FE89",
X"FE89",
X"FE0C",
X"FF06",
X"FF06",
X"0000",
X"00FA",
X"007D",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"007D",
X"00FA",
X"01F4",
X"02EE",
X"036B",
X"02EE",
X"02EE",
X"0465",
X"0465",
X"03E8",
X"0465",
X"05DC",
X"055F",
X"0465",
X"055F",
X"055F",
X"03E8",
X"055F",
X"0659",
X"055F",
X"03E8",
X"055F",
X"04E2",
X"03E8",
X"04E2",
X"04E2",
X"055F",
X"0465",
X"036B",
X"0465",
X"03E8",
X"03E8",
X"03E8",
X"0465",
X"0465",
X"0465",
X"0465",
X"055F",
X"055F",
X"05DC",
X"06D6",
X"05DC",
X"06D6",
X"06D6",
X"06D6",
X"0659",
X"06D6",
X"0753",
X"0659",
X"06D6",
X"0659",
X"05DC",
X"055F",
X"05DC",
X"05DC",
X"0465",
X"05DC",
X"0659",
X"0659",
X"0659",
X"0659",
X"06D6",
X"06D6",
X"06D6",
X"0659",
X"0753",
X"06D6",
X"06D6",
X"06D6",
X"06D6",
X"06D6",
X"0659",
X"06D6",
X"0659",
X"0659",
X"0659",
X"0659",
X"055F",
X"04E2",
X"03E8",
X"036B",
X"036B",
X"03E8",
X"036B",
X"036B",
X"036B",
X"036B",
X"02EE",
X"02EE",
X"0271",
X"0177",
X"00FA",
X"0177",
X"007D",
X"FF83",
X"00FA",
X"007D",
X"FF83",
X"FF83",
X"FF83",
X"FE89",
X"FC18",
X"FC95",
X"FB1E",
X"FB1E",
X"FB1E",
X"FAA1",
X"FB1E",
X"FB1E",
X"FA24",
X"FB1E",
X"FA24",
X"FA24",
X"F9A7",
X"F92A",
X"FA24",
X"F92A",
X"F92A",
X"FA24",
X"F9A7",
X"F9A7",
X"F9A7",
X"FA24",
X"FA24",
X"F8AD",
X"F92A",
X"FA24",
X"F9A7",
X"F9A7",
X"F8AD",
X"F92A",
X"FA24",
X"FA24",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB9B",
X"FB9B",
X"FB9B",
X"FC18",
X"FB9B",
X"FD12",
X"FC95",
X"FC18",
X"FD8F",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FB9B",
X"FB1E",
X"FB1E",
X"FAA1",
X"FAA1",
X"FB9B",
X"FB1E",
X"FA24",
X"FA24",
X"FAA1",
X"FAA1",
X"FA24",
X"F9A7",
X"F8AD",
X"F92A",
X"F9A7",
X"FA24",
X"F9A7",
X"FA24",
X"F9A7",
X"FA24",
X"FB1E",
X"FA24",
X"FAA1",
X"FB1E",
X"FB1E",
X"FA24",
X"F9A7",
X"FA24",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FD12",
X"FE0C",
X"FE89",
X"FF83",
X"0000",
X"007D",
X"007D",
X"0177",
X"01F4",
X"01F4",
X"0177",
X"0271",
X"0271",
X"01F4",
X"02EE",
X"02EE",
X"03E8",
X"03E8",
X"036B",
X"03E8",
X"0465",
X"04E2",
X"0465",
X"04E2",
X"055F",
X"04E2",
X"04E2",
X"05DC",
X"05DC",
X"0465",
X"0465",
X"04E2",
X"0465",
X"055F",
X"04E2",
X"03E8",
X"04E2",
X"055F",
X"055F",
X"04E2",
X"0465",
X"036B",
X"036B",
X"0271",
X"0271",
X"0271",
X"0271",
X"02EE",
X"0271",
X"02EE",
X"036B",
X"036B",
X"02EE",
X"036B",
X"02EE",
X"01F4",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"0000",
X"00FA",
X"FF83",
X"FF06",
X"00FA",
X"00FA",
X"FF06",
X"FE89",
X"0000",
X"FF06",
X"FE89",
X"FE89",
X"FE0C",
X"FD8F",
X"FE89",
X"FE0C",
X"FF06",
X"FF83",
X"FF06",
X"FF83",
X"FF06",
X"0000",
X"007D",
X"007D",
X"FF06",
X"FF83",
X"0000",
X"FF83",
X"0000",
X"007D",
X"0177",
X"01F4",
X"0177",
X"00FA",
X"01F4",
X"01F4",
X"00FA",
X"01F4",
X"01F4",
X"01F4",
X"03E8",
X"02EE",
X"01F4",
X"0271",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"036B",
X"03E8",
X"02EE",
X"0271",
X"02EE",
X"0271",
X"0177",
X"01F4",
X"0271",
X"0271",
X"0271",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"02EE",
X"02EE",
X"0271",
X"02EE",
X"02EE",
X"0271",
X"0271",
X"02EE",
X"01F4",
X"01F4",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"0271",
X"0271",
X"036B",
X"0271",
X"01F4",
X"0271",
X"02EE",
X"02EE",
X"0271",
X"00FA",
X"0177",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"00FA",
X"007D",
X"007D",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FD12",
X"FD8F",
X"FE89",
X"FD12",
X"FC95",
X"FC18",
X"FC95",
X"FC95",
X"FD12",
X"FC18",
X"FC95",
X"FD8F",
X"FC95",
X"FC18",
X"FC95",
X"FD12",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FE0C",
X"FD8F",
X"FD12",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE0C",
X"FD8F",
X"FF06",
X"0000",
X"FE89",
X"FE0C",
X"007D",
X"0000",
X"FD8F",
X"FE89",
X"FF83",
X"FF83",
X"FE0C",
X"FD8F",
X"FE89",
X"FE89",
X"FE0C",
X"FD12",
X"FE89",
X"FF06",
X"FE89",
X"FD8F",
X"FE89",
X"FF06",
X"FD12",
X"FD8F",
X"FF83",
X"FE0C",
X"FC95",
X"FE0C",
X"FD12",
X"FC18",
X"FB9B",
X"FC95",
X"FD8F",
X"FC95",
X"FC18",
X"FC95",
X"FB9B",
X"FB1E",
X"FC18",
X"FC18",
X"FAA1",
X"FC18",
X"FC95",
X"FC95",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE89",
X"FE0C",
X"FF83",
X"0000",
X"FF06",
X"0000",
X"0000",
X"FF83",
X"0000",
X"FF83",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"00FA",
X"01F4",
X"0271",
X"01F4",
X"01F4",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"036B",
X"0271",
X"01F4",
X"02EE",
X"02EE",
X"0271",
X"0271",
X"01F4",
X"02EE",
X"0271",
X"01F4",
X"02EE",
X"02EE",
X"01F4",
X"0177",
X"01F4",
X"0177",
X"0271",
X"0177",
X"00FA",
X"01F4",
X"0271",
X"01F4",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"00FA",
X"01F4",
X"0271",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"007D",
X"007D",
X"007D",
X"FF83",
X"FF83",
X"0000",
X"FE89",
X"FE89",
X"FE89",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD12",
X"FD8F",
X"FD8F",
X"FD12",
X"FD8F",
X"FE0C",
X"FD8F",
X"FD12",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC95",
X"FC18",
X"FC95",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE89",
X"FE0C",
X"FE0C",
X"FD8F",
X"FE89",
X"FF83",
X"FF06",
X"FE89",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF83",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"007D",
X"0000",
X"0000",
X"007D",
X"0000",
X"007D",
X"007D",
X"007D",
X"0177",
X"0177",
X"0177",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"03E8",
X"0465",
X"0465",
X"03E8",
X"0465",
X"04E2",
X"04E2",
X"0465",
X"0465",
X"0465",
X"04E2",
X"055F",
X"04E2",
X"055F",
X"0659",
X"06D6",
X"07D0",
X"07D0",
X"0753",
X"0753",
X"06D6",
X"0659",
X"0753",
X"0753",
X"0753",
X"06D6",
X"0659",
X"06D6",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"04E2",
X"055F",
X"055F",
X"04E2",
X"04E2",
X"055F",
X"055F",
X"0465",
X"036B",
X"036B",
X"02EE",
X"0271",
X"0271",
X"0271",
X"01F4",
X"0177",
X"00FA",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"FD8F",
X"FE0C",
X"FE0C",
X"FC18",
X"FC95",
X"FD12",
X"FD12",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FB9B",
X"FAA1",
X"FAA1",
X"FAA1",
X"FAA1",
X"FA24",
X"FA24",
X"FA24",
X"FAA1",
X"FA24",
X"FA24",
X"FAA1",
X"FAA1",
X"FAA1",
X"FB1E",
X"FAA1",
X"FA24",
X"F9A7",
X"F9A7",
X"F92A",
X"F92A",
X"FA24",
X"F92A",
X"F9A7",
X"FB9B",
X"FAA1",
X"FB1E",
X"FC18",
X"FC95",
X"FC95",
X"FC95",
X"FB9B",
X"FA24",
X"FB1E",
X"FB9B",
X"FC18",
X"FAA1",
X"F9A7",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FB1E",
X"FC95",
X"FD8F",
X"FC95",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FD8F",
X"FF83",
X"FE89",
X"FE89",
X"FF83",
X"FF06",
X"FE89",
X"FF83",
X"FF83",
X"007D",
X"0000",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"01F4",
X"0177",
X"007D",
X"01F4",
X"01F4",
X"0177",
X"0271",
X"01F4",
X"00FA",
X"00FA",
X"0177",
X"00FA",
X"0000",
X"007D",
X"007D",
X"007D",
X"00FA",
X"0177",
X"007D",
X"007D",
X"00FA",
X"007D",
X"FF83",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"01F4",
X"0000",
X"007D",
X"0177",
X"007D",
X"00FA",
X"007D",
X"00FA",
X"00FA",
X"007D",
X"00FA",
X"007D",
X"007D",
X"007D",
X"00FA",
X"0000",
X"0000",
X"007D",
X"00FA",
X"007D",
X"0000",
X"007D",
X"007D",
X"FF83",
X"007D",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"007D",
X"0177",
X"0177",
X"007D",
X"00FA",
X"01F4",
X"01F4",
X"0271",
X"036B",
X"02EE",
X"02EE",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"02EE",
X"036B",
X"0271",
X"036B",
X"03E8",
X"03E8",
X"036B",
X"036B",
X"036B",
X"03E8",
X"0465",
X"036B",
X"0465",
X"036B",
X"03E8",
X"03E8",
X"0271",
X"0271",
X"01F4",
X"0177",
X"0177",
X"007D",
X"00FA",
X"0000",
X"007D",
X"00FA",
X"FF83",
X"FF83",
X"FF06",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FE0C",
X"FF83",
X"FF83",
X"FE89",
X"FF06",
X"FF83",
X"FF06",
X"FE89",
X"FF06",
X"FF06",
X"FE89",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FE89",
X"FE0C",
X"FE89",
X"FF06",
X"FE89",
X"FF06",
X"FE89",
X"FE89",
X"FE0C",
X"FD8F",
X"FD12",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FC95",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FE0C",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FD8F",
X"FE0C",
X"FE89",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"FF83",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"FF83",
X"0000",
X"007D",
X"007D",
X"0000",
X"007D",
X"00FA",
X"0177",
X"0177",
X"01F4",
X"0271",
X"0271",
X"0271",
X"0271",
X"02EE",
X"0271",
X"0271",
X"02EE",
X"0271",
X"0271",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"0271",
X"02EE",
X"036B",
X"036B",
X"036B",
X"02EE",
X"02EE",
X"036B",
X"02EE",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"02EE",
X"0271",
X"02EE",
X"0271",
X"01F4",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF06",
X"FF83",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"FF83",
X"0000",
X"007D",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0271",
X"02EE",
X"0271",
X"02EE",
X"0271",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"02EE",
X"0271",
X"0271",
X"02EE",
X"02EE",
X"01F4",
X"01F4",
X"0177",
X"01F4",
X"01F4",
X"0177",
X"00FA",
X"00FA",
X"0177",
X"007D",
X"0000",
X"0000",
X"007D",
X"0000",
X"FF83",
X"0000",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD12",
X"FC18",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF83",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FE89",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD8F",
X"FD12",
X"FC18",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FB1E",
X"FB9B",
X"FB9B",
X"FB1E",
X"FC18",
X"FC18",
X"FC95",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"0271",
X"01F4",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"0271",
X"02EE",
X"036B",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"03E8",
X"0465",
X"0465",
X"0465",
X"04E2",
X"04E2",
X"04E2",
X"055F",
X"055F",
X"05DC",
X"05DC",
X"05DC",
X"0659",
X"06D6",
X"0659",
X"0659",
X"05DC",
X"05DC",
X"0659",
X"05DC",
X"05DC",
X"055F",
X"0465",
X"04E2",
X"0465",
X"03E8",
X"0465",
X"0465",
X"03E8",
X"03E8",
X"036B",
X"02EE",
X"02EE",
X"036B",
X"02EE",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"0271",
X"01F4",
X"0271",
X"0271",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0271",
X"02EE",
X"02EE",
X"036B",
X"036B",
X"03E8",
X"03E8",
X"03E8",
X"036B",
X"036B",
X"0465",
X"036B",
X"02EE",
X"02EE",
X"02EE",
X"0271",
X"0177",
X"0177",
X"01F4",
X"0177",
X"0177",
X"00FA",
X"007D",
X"00FA",
X"007D",
X"00FA",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FE89",
X"FE89",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD12",
X"FC95",
X"FD12",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC95",
X"FC18",
X"FC18",
X"FC18",
X"FB9B",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB1E",
X"FB9B",
X"FB1E",
X"FB9B",
X"FB9B",
X"FB1E",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FB9B",
X"FC18",
X"FB9B",
X"FC18",
X"FC18",
X"FC18",
X"FC18",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FC95",
X"FD12",
X"FC95",
X"FD12",
X"FD8F",
X"FD12",
X"FD8F",
X"FC95",
X"FD12",
X"FD8F",
X"FE0C",
X"FD8F",
X"FD12",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD8F",
X"FE0C",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD12",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD12",
X"FD8F",
X"FC95",
X"FD12",
X"FD8F",
X"FD8F",
X"FE0C",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE89",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"FF06",
X"FE89",
X"FF83",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"0177",
X"00FA",
X"0177",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"0271",
X"0271",
X"02EE",
X"036B",
X"03E8",
X"036B",
X"036B",
X"03E8",
X"0465",
X"0465",
X"03E8",
X"03E8",
X"03E8",
X"0465",
X"0465",
X"04E2",
X"0465",
X"0465",
X"04E2",
X"055F",
X"055F",
X"055F",
X"04E2",
X"055F",
X"05DC",
X"05DC",
X"05DC",
X"05DC",
X"0659",
X"05DC",
X"0659",
X"0659",
X"05DC",
X"05DC",
X"05DC",
X"055F",
X"05DC",
X"0659",
X"05DC",
X"0659",
X"05DC",
X"05DC",
X"04E2",
X"04E2",
X"055F",
X"04E2",
X"03E8",
X"036B",
X"036B",
X"03E8",
X"036B",
X"02EE",
X"036B",
X"02EE",
X"0271",
X"02EE",
X"02EE",
X"02EE",
X"0271",
X"0271",
X"0271",
X"0271",
X"01F4",
X"0271",
X"01F4",
X"0271",
X"01F4",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"007D",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"FF83",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF06",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE0C",
X"FD8F",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FC18",
X"FC95",
X"FC18",
X"FC95",
X"FD12",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FC95",
X"FC18",
X"FC18",
X"FC95",
X"FC18",
X"FC18",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FC95",
X"FD12",
X"FD12",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FC95",
X"FC95",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD12",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FC95",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FE0C",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE0C",
X"FF06",
X"FE89",
X"FE0C",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"0000",
X"0000",
X"FF83",
X"00FA",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"0177",
X"01F4",
X"0177",
X"01F4",
X"0271",
X"0271",
X"02EE",
X"02EE",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"036B",
X"02EE",
X"02EE",
X"036B",
X"036B",
X"02EE",
X"02EE",
X"036B",
X"036B",
X"036B",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"02EE",
X"0271",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"01F4",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"01F4",
X"0177",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"00FA",
X"0177",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"007D",
X"007D",
X"0000",
X"007D",
X"007D",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FD8F",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF83",
X"FE89",
X"FF06",
X"FE89",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"FF83",
X"0000",
X"0000",
X"FF06",
X"FF06",
X"0000",
X"FF06",
X"FE89",
X"FF83",
X"FF83",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF83",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"01F4",
X"0271",
X"0177",
X"0177",
X"0271",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"0271",
X"02EE",
X"02EE",
X"0271",
X"01F4",
X"0271",
X"01F4",
X"0271",
X"01F4",
X"0177",
X"00FA",
X"01F4",
X"01F4",
X"00FA",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"0177",
X"00FA",
X"00FA",
X"0000",
X"0000",
X"007D",
X"0000",
X"007D",
X"00FA",
X"0177",
X"0177",
X"01F4",
X"0177",
X"0177",
X"01F4",
X"00FA",
X"0177",
X"007D",
X"FF06",
X"FF83",
X"007D",
X"007D",
X"0000",
X"007D",
X"00FA",
X"007D",
X"FF83",
X"FF83",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FF83",
X"FF06",
X"FF83",
X"FF83",
X"FF06",
X"FE89",
X"FE89",
X"FF06",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FE89",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"FF06",
X"FF83",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"0000",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"01F4",
X"0177",
X"0177",
X"0177",
X"0177",
X"01F4",
X"0177",
X"0177",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0000",
X"007D",
X"0000",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD8F",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD12",
X"FD8F",
X"FD12",
X"FD8F",
X"FD8F",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"007D",
X"00FA",
X"0177",
X"01F4",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"00FA",
X"007D",
X"007D",
X"007D",
X"00FA",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"0000",
X"007D",
X"0000",
X"0000",
X"0000",
X"FF06",
X"0000",
X"0000",
X"0000",
X"FF83",
X"0000",
X"007D",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"00FA",
X"0177",
X"00FA",
X"00FA",
X"0000",
X"0177",
X"01F4",
X"0177",
X"0177",
X"00FA",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"0271",
X"02EE",
X"00FA",
X"00FA",
X"01F4",
X"0271",
X"01F4",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"0000",
X"0000",
X"00FA",
X"0177",
X"007D",
X"0000",
X"007D",
X"007D",
X"007D",
X"00FA",
X"FF83",
X"FF83",
X"007D",
X"00FA",
X"0000",
X"FF83",
X"0000",
X"FF06",
X"FF06",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FE89",
X"FE0C",
X"FE89",
X"FF83",
X"FF06",
X"FD8F",
X"FD8F",
X"FE89",
X"FF06",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FE0C",
X"FD8F",
X"FD8F",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FE0C",
X"FE89",
X"FF06",
X"FF06",
X"FF06",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FF06",
X"FE89",
X"FE0C",
X"FE0C",
X"FF06",
X"FF83",
X"FF83",
X"FE89",
X"FE89",
X"FF83",
X"FF06",
X"FF83",
X"0000",
X"0000",
X"FF83",
X"0000",
X"FF06",
X"FE89",
X"FF06",
X"FF83",
X"FF83",
X"FE89",
X"FF83",
X"FF83",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF06",
X"007D",
X"0000",
X"FE89",
X"FE89",
X"FF83",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"FF83",
X"FF06",
X"0000",
X"0000",
X"FF83",
X"0000",
X"00FA",
X"007D",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"007D",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"0000",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"0000",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"0177",
X"01F4",
X"0177",
X"007D",
X"00FA",
X"01F4",
X"01F4",
X"0177",
X"01F4",
X"0271",
X"0271",
X"01F4",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"01F4",
X"0271",
X"0271",
X"0271",
X"0271",
X"0177",
X"01F4",
X"0271",
X"01F4",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"0177",
X"01F4",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"00FA",
X"007D",
X"007D",
X"007D",
X"0177",
X"00FA",
X"007D",
X"007D",
X"00FA",
X"007D",
X"007D",
X"007D",
X"0000",
X"FF83",
X"007D",
X"007D",
X"FF06",
X"0000",
X"0000",
X"FF06",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"00FA",
X"007D",
X"FE89",
X"FF06",
X"0000",
X"007D",
X"FF83",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"FE89",
X"FF83",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FF83",
X"FF83",
X"FF06",
X"0000",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FE89",
X"FF06",
X"FF83",
X"FE89",
X"FE0C",
X"FE0C",
X"FF06",
X"0000",
X"0000",
X"FF06",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"0000",
X"FF83",
X"FE89",
X"FE89",
X"FF06",
X"FF83",
X"FF06",
X"FE89",
X"FF06",
X"0000",
X"0000",
X"FF06",
X"FF83",
X"0000",
X"FF83",
X"0000",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"007D",
X"00FA",
X"0000",
X"0000",
X"FF06",
X"FF83",
X"007D",
X"007D",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"0000",
X"FF83",
X"FE89",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FE89",
X"FE0C",
X"FE89",
X"FF06",
X"FF83",
X"FE0C",
X"FE0C",
X"FE89",
X"FF06",
X"FE89",
X"FD8F",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF83",
X"FE89",
X"FE89",
X"0000",
X"0000",
X"FF83",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"FF83",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"FF06",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"0000",
X"FF83",
X"FF06",
X"FF83",
X"007D",
X"007D",
X"FF83",
X"FF06",
X"FF83",
X"007D",
X"007D",
X"FF83",
X"FF83",
X"007D",
X"007D",
X"FF83",
X"007D",
X"0000",
X"0000",
X"00FA",
X"007D",
X"0000",
X"00FA",
X"00FA",
X"0000",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"00FA",
X"007D",
X"01F4",
X"01F4",
X"0177",
X"00FA",
X"0000",
X"007D",
X"0177",
X"0177",
X"0177",
X"007D",
X"00FA",
X"01F4",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"0177",
X"00FA",
X"0177",
X"00FA",
X"0177",
X"0177",
X"00FA",
X"0177",
X"00FA",
X"007D",
X"00FA",
X"00FA",
X"007D",
X"00FA",
X"0000",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"0000",
X"FF83",
X"007D",
X"00FA",
X"007D",
X"FF83",
X"FF83",
X"0000",
X"007D",
X"00FA",
X"0000",
X"0000",
X"007D",
X"007D",
X"0000",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"00FA",
X"0177",
X"0177",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"0177",
X"00FA",
X"0177",
X"00FA",
X"007D",
X"00FA",
X"01F4",
X"0271",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"00FA",
X"01F4",
X"0177",
X"007D",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FE89",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF06",
X"FF83",
X"0000",
X"FF83",
X"FF06",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF83",
X"FF06",
X"FF06",
X"FF83",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE0C",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE0C",
X"FF06",
X"FF06",
X"FE0C",
X"FE89",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"0000",
X"FF83",
X"FF06",
X"0000",
X"0000",
X"FF83",
X"0000",
X"0000",
X"0000",
X"FF83",
X"0000",
X"007D",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"00FA",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"01F4",
X"0177",
X"0177",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"0271",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"0271",
X"01F4",
X"0271",
X"0271",
X"01F4",
X"0271",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"01F4",
X"0177",
X"01F4",
X"01F4",
X"0177",
X"0177",
X"0177",
X"01F4",
X"0177",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FE89",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE0C",
X"FE0C",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FE89",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"007D",
X"007D",
X"0000",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"FF83",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"0000",
X"007D",
X"0000",
X"0000",
X"007D",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"007D",
X"007D",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"01F4",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"00FA",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"0177",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"00FA",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FE89",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"FF83",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"00FA",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"00FA",
X"00FA",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"007D",
X"007D",
X"0000",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"0000",
X"0000",
X"FF83",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE0C",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"0177",
X"00FA",
X"00FA",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"0177",
X"00FA",
X"0177",
X"0177",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FE89",
X"FF06",
X"FE89",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"FF83",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"00FA",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"00FA",
X"00FA",
X"007D",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"0000",
X"0000",
X"007D",
X"007D",
X"0000",
X"007D",
X"007D",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"0000",
X"0000",
X"FF83",
X"0000",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"FF83",
X"FF83",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF06",
X"FF06",
X"FF83",
X"FF06",
X"FF06",
X"FF06",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"FF83",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"007D",
X"0000",
X"0000",
X"0000",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"00FA",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D",
X"007D"





 );

 
 begin

    if (resetN='0') then
		Q_tmp <= ( others => '0');
    elsif(rising_edge(CLK)) then
      if (ENA='1') then
		Q_tmp <= sin_table(conv_integer(ADDR));
		else 
	 Q_tmp <= ( others => '0');
      end if;
   end if;
  end process;
 Q <= Q_tmp; 

		   
end arch;