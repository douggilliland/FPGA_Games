-- generated with romgen v3.03 by MikeJ
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_unsigned.all;
	use ieee.numeric_std.all;

library UNISIM;
	use UNISIM.Vcomponents.all;

entity ROM_D2 is
port (
	CLK  : in  std_logic;
	ADDR : in  std_logic_vector(10 downto 0);
	DATA : out std_logic_vector(7 downto 0)
	);
end;

architecture RTL of ROM_D2 is


	type ROM_ARRAY is array(0 to 2047) of std_logic_vector(7 downto 0);
	constant ROM : ROM_ARRAY := (
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0000
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0008
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0010
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0018
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0020
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0028
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0030
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0038
		x"40",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0040
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0048
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0050
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0058
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0060
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0068
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0070
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0078
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0080
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0088
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0090
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"01", -- 0x0098
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x00A0
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x00A8
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x00B0
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"1E", -- 0x00B8
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x00C0
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x00C8
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x00D0
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"19", -- 0x00D8
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x00E0
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x00E8
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x00F0
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x00F8
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0100
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0108
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0110
		x"30",x"30",x"30",x"30",x"30",x"30",x"00",x"30", -- 0x0118
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0120
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0128
		x"30",x"15",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0130
		x"30",x"30",x"30",x"30",x"30",x"30",x"00",x"30", -- 0x0138
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0140
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0148
		x"30",x"0A",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0150
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0158
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0160
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0168
		x"30",x"1C",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0170
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"11", -- 0x0178
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0180
		x"30",x"30",x"30",x"19",x"30",x"30",x"30",x"30", -- 0x0188
		x"30",x"1D",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0190
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"12", -- 0x0198
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x01A0
		x"30",x"30",x"30",x"15",x"30",x"1B",x"30",x"30", -- 0x01A8
		x"30",x"30",x"30",x"30",x"16",x"30",x"30",x"30", -- 0x01B0
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"10", -- 0x01B8
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x01C0
		x"30",x"30",x"30",x"0A",x"30",x"0E",x"30",x"30", -- 0x01C8
		x"30",x"03",x"30",x"30",x"12",x"30",x"30",x"30", -- 0x01D0
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"11", -- 0x01D8
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x01E0
		x"30",x"30",x"30",x"22",x"30",x"0A",x"30",x"30", -- 0x01E8
		x"30",x"02",x"30",x"30",x"0D",x"30",x"30",x"30", -- 0x01F0
		x"30",x"30",x"30",x"30",x"30",x"30",x"04",x"30", -- 0x01F8
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0200
		x"30",x"30",x"30",x"0E",x"30",x"0D",x"30",x"30", -- 0x0208
		x"30",x"30",x"30",x"30",x"20",x"30",x"30",x"30", -- 0x0210
		x"30",x"30",x"30",x"30",x"30",x"30",x"00",x"1C", -- 0x0218
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0220
		x"30",x"30",x"30",x"1B",x"30",x"22",x"30",x"30", -- 0x0228
		x"30",x"1C",x"30",x"30",x"0A",x"30",x"30",x"30", -- 0x0230
		x"30",x"30",x"30",x"30",x"30",x"30",x"00",x"0C", -- 0x0238
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0240
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0248
		x"30",x"1D",x"30",x"30",x"22",x"30",x"30",x"30", -- 0x0250
		x"30",x"30",x"30",x"30",x"30",x"30",x"00",x"18", -- 0x0258
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0260
		x"30",x"30",x"30",x"01",x"30",x"30",x"30",x"30", -- 0x0268
		x"30",x"0A",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0270
		x"30",x"30",x"30",x"30",x"30",x"30",x"00",x"1B", -- 0x0278
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0280
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0288
		x"30",x"10",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0290
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"0E", -- 0x0298
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x02A0
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x02A8
		x"30",x"0E",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x02B0
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x02B8
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x02C0
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x02C8
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x02D0
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x02D8
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x02E0
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x02E8
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x02F0
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x02F8
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0300
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0308
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0310
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0318
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0320
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0328
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0330
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"02", -- 0x0338
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0340
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0348
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0350
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"1E", -- 0x0358
		x"68",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0360
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0368
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0370
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"19", -- 0x0378
		x"68",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0380
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0388
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0390
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x0398
		x"68",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x03A0
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x03A8
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x03B0
		x"30",x"30",x"30",x"30",x"30",x"30",x"30",x"30", -- 0x03B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x03F8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0400
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0408
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0410
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0418
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0420
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0428
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0430
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0438
		x"32",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0440
		x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C", -- 0x0448
		x"00",x"1A",x"00",x"00",x"16",x"00",x"00",x"00", -- 0x0450
		x"00",x"19",x"00",x"00",x"00",x"00",x"33",x"19", -- 0x0458
		x"32",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0460
		x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C", -- 0x0468
		x"00",x"1A",x"00",x"00",x"16",x"00",x"00",x"00", -- 0x0470
		x"00",x"19",x"00",x"00",x"00",x"00",x"33",x"19", -- 0x0478
		x"32",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0480
		x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C", -- 0x0488
		x"00",x"1A",x"00",x"00",x"16",x"00",x"00",x"00", -- 0x0490
		x"00",x"19",x"00",x"00",x"00",x"00",x"33",x"19", -- 0x0498
		x"32",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04A0
		x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C", -- 0x04A8
		x"00",x"1A",x"00",x"00",x"16",x"00",x"00",x"00", -- 0x04B0
		x"00",x"19",x"00",x"00",x"00",x"00",x"33",x"19", -- 0x04B8
		x"32",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04C0
		x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C", -- 0x04C8
		x"00",x"1A",x"00",x"00",x"16",x"00",x"00",x"00", -- 0x04D0
		x"00",x"19",x"00",x"00",x"00",x"00",x"33",x"19", -- 0x04D8
		x"32",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x04E0
		x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C", -- 0x04E8
		x"00",x"1A",x"00",x"00",x"16",x"00",x"00",x"00", -- 0x04F0
		x"00",x"19",x"00",x"00",x"00",x"00",x"33",x"19", -- 0x04F8
		x"32",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0500
		x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C", -- 0x0508
		x"00",x"1A",x"00",x"00",x"16",x"00",x"00",x"00", -- 0x0510
		x"00",x"19",x"00",x"00",x"00",x"00",x"33",x"19", -- 0x0518
		x"32",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0520
		x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C", -- 0x0528
		x"00",x"1A",x"00",x"00",x"16",x"00",x"00",x"00", -- 0x0530
		x"00",x"19",x"00",x"00",x"00",x"00",x"33",x"19", -- 0x0538
		x"32",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0540
		x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C", -- 0x0548
		x"00",x"1A",x"00",x"00",x"16",x"00",x"00",x"00", -- 0x0550
		x"00",x"19",x"00",x"00",x"00",x"00",x"33",x"19", -- 0x0558
		x"32",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0560
		x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C", -- 0x0568
		x"00",x"1A",x"00",x"00",x"16",x"00",x"00",x"00", -- 0x0570
		x"00",x"19",x"00",x"00",x"00",x"00",x"33",x"1A", -- 0x0578
		x"32",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0580
		x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C", -- 0x0588
		x"00",x"1A",x"00",x"00",x"16",x"00",x"00",x"00", -- 0x0590
		x"00",x"19",x"00",x"00",x"00",x"00",x"33",x"1A", -- 0x0598
		x"32",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05A0
		x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C", -- 0x05A8
		x"00",x"1A",x"00",x"00",x"16",x"00",x"00",x"00", -- 0x05B0
		x"00",x"19",x"00",x"00",x"00",x"00",x"33",x"1A", -- 0x05B8
		x"32",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05C0
		x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C", -- 0x05C8
		x"00",x"1A",x"00",x"00",x"16",x"00",x"00",x"00", -- 0x05D0
		x"00",x"19",x"00",x"00",x"00",x"00",x"33",x"1A", -- 0x05D8
		x"32",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x05E0
		x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C", -- 0x05E8
		x"00",x"1A",x"00",x"00",x"16",x"00",x"00",x"00", -- 0x05F0
		x"00",x"19",x"00",x"00",x"00",x"00",x"33",x"1A", -- 0x05F8
		x"32",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0600
		x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C", -- 0x0608
		x"00",x"1A",x"00",x"00",x"16",x"00",x"00",x"00", -- 0x0610
		x"00",x"19",x"00",x"00",x"00",x"00",x"33",x"1A", -- 0x0618
		x"32",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0620
		x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C", -- 0x0628
		x"00",x"1A",x"00",x"00",x"16",x"00",x"00",x"00", -- 0x0630
		x"00",x"19",x"00",x"00",x"00",x"00",x"33",x"1A", -- 0x0638
		x"32",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0640
		x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C", -- 0x0648
		x"00",x"1A",x"00",x"00",x"16",x"00",x"00",x"00", -- 0x0650
		x"00",x"19",x"00",x"00",x"00",x"00",x"33",x"1A", -- 0x0658
		x"32",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0660
		x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C", -- 0x0668
		x"00",x"1A",x"00",x"00",x"16",x"00",x"00",x"00", -- 0x0670
		x"00",x"19",x"00",x"00",x"00",x"00",x"33",x"1A", -- 0x0678
		x"32",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0680
		x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C", -- 0x0688
		x"00",x"1A",x"00",x"00",x"16",x"00",x"00",x"00", -- 0x0690
		x"00",x"19",x"00",x"00",x"00",x"00",x"33",x"1A", -- 0x0698
		x"32",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06A0
		x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C", -- 0x06A8
		x"00",x"1A",x"00",x"00",x"16",x"00",x"00",x"00", -- 0x06B0
		x"00",x"19",x"00",x"00",x"00",x"00",x"33",x"19", -- 0x06B8
		x"32",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06C0
		x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C", -- 0x06C8
		x"00",x"1A",x"00",x"00",x"16",x"00",x"00",x"00", -- 0x06D0
		x"00",x"19",x"00",x"00",x"00",x"00",x"33",x"19", -- 0x06D8
		x"32",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x06E0
		x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C", -- 0x06E8
		x"00",x"1A",x"00",x"00",x"16",x"00",x"00",x"00", -- 0x06F0
		x"00",x"19",x"00",x"00",x"00",x"00",x"33",x"19", -- 0x06F8
		x"05",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0700
		x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C", -- 0x0708
		x"00",x"1A",x"00",x"00",x"16",x"00",x"00",x"00", -- 0x0710
		x"00",x"19",x"00",x"00",x"00",x"00",x"33",x"19", -- 0x0718
		x"05",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0720
		x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C", -- 0x0728
		x"00",x"1A",x"00",x"00",x"16",x"00",x"00",x"00", -- 0x0730
		x"00",x"19",x"00",x"00",x"00",x"00",x"33",x"00", -- 0x0738
		x"05",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0740
		x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C", -- 0x0748
		x"00",x"1A",x"00",x"00",x"16",x"00",x"00",x"00", -- 0x0750
		x"00",x"19",x"00",x"00",x"00",x"00",x"33",x"00", -- 0x0758
		x"05",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0760
		x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C", -- 0x0768
		x"00",x"1A",x"00",x"00",x"16",x"00",x"00",x"00", -- 0x0770
		x"00",x"19",x"00",x"00",x"00",x"00",x"33",x"00", -- 0x0778
		x"05",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x0780
		x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C", -- 0x0788
		x"00",x"1A",x"00",x"00",x"16",x"00",x"00",x"00", -- 0x0790
		x"00",x"19",x"00",x"00",x"00",x"00",x"33",x"19", -- 0x0798
		x"05",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07A0
		x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C",x"3C", -- 0x07A8
		x"00",x"1A",x"00",x"00",x"16",x"00",x"00",x"00", -- 0x07B0
		x"00",x"19",x"00",x"00",x"00",x"00",x"33",x"19", -- 0x07B8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07C0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07C8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07D0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07D8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07E0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07E8
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 0x07F0
		x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00"  -- 0x07F8
	);

begin

	p_rom : process
	begin
		wait until rising_edge(CLK);
			DATA <= ROM(to_integer(unsigned(ADDR)));
	end process;
end RTL;
