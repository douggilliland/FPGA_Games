library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


entity Car1_drawer is 
	Port(
		 
		 DrawX: in std_logic_vector( 9 downto 0); 
		 DrawY: in std_logic_vector( 9 downto 0);
		 Car_X_center: in std_logic_vector (9 downto 0); 
		 Car_Y_center: in std_logic_vector (9 downto 0); 
		 draw_red: out std_logic_vector(7 downto 0);
		 draw_green: out std_logic_vector(7 downto 0);
		 draw_blue: out std_logic_vector(7 downto 0)
		 
		 );
end entity;



architecture table of Car1_drawer is

type car is array (1199 downto 0) of std_logic_vector(7 downto 0);
signal car_red : car := (

x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"05",
x"01",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"0f",
x"03",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"0c",
x"0f",
x"0f",
x"0f",
x"0f",
x"0f",
x"06",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"02",
x"0f",
x"0f",
x"0f",
x"0f",
x"0f",
x"02",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"0d",
x"5b",
x"7d",
x"7e",
x"7e",
x"7e",
x"75",
x"40",
x"09",
x"10",
x"01",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"0c",
x"62",
x"77",
x"75",
x"7e",
x"71",
x"31",
x"02",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"20",
x"36",
x"24",
x"76",
x"a7",
x"a9",
x"a9",
x"a9",
x"99",
x"5c",
x"32",
x"5c",
x"5b",
x"5a",
x"5a",
x"5a",
x"5a",
x"5a",
x"36",
x"05",
x"25",
x"8a",
x"9d",
x"8e",
x"ae",
x"d9",
x"93",
x"2e",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"09",
x"54",
x"82",
x"3a",
x"2e",
x"36",
x"3b",
x"51",
x"46",
x"34",
x"2a",
x"4d",
x"a8",
x"b5",
x"b5",
x"b5",
x"b5",
x"b5",
x"b5",
x"6d",
x"21",
x"3d",
x"46",
x"3e",
x"3e",
x"58",
x"b2",
x"bd",
x"5a",
x"15",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"06",
x"13",
x"16",
x"3e",
x"45",
x"44",
x"29",
x"2c",
x"44",
x"34",
x"25",
x"16",
x"23",
x"61",
x"4b",
x"2c",
x"28",
x"29",
x"28",
x"3b",
x"2b",
x"20",
x"24",
x"23",
x"37",
x"4c",
x"3f",
x"44",
x"4c",
x"0e",
x"02",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"02",
x"42",
x"95",
x"a0",
x"a0",
x"a0",
x"a5",
x"85",
x"40",
x"71",
x"a4",
x"a6",
x"a6",
x"9b",
x"54",
x"15",
x"1e",
x"0c",
x"00",
x"19",
x"21",
x"3a",
x"3a",
x"2e",
x"2a",
x"2b",
x"24",
x"87",
x"5c",
x"05",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"08",
x"4a",
x"84",
x"7d",
x"7a",
x"7b",
x"8d",
x"67",
x"37",
x"5e",
x"8c",
x"98",
x"9a",
x"84",
x"7f",
x"61",
x"1b",
x"09",
x"03",
x"12",
x"1f",
x"1f",
x"19",
x"14",
x"10",
x"20",
x"29",
x"5b",
x"42",
x"12",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"18",
x"33",
x"2f",
x"22",
x"2c",
x"20",
x"20",
x"20",
x"30",
x"2c",
x"2e",
x"3e",
x"3a",
x"8d",
x"96",
x"2c",
x"13",
x"06",
x"2a",
x"52",
x"52",
x"47",
x"4e",
x"4b",
x"5d",
x"4b",
x"52",
x"26",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"04",
x"0b",
x"0f",
x"20",
x"2a",
x"23",
x"2d",
x"20",
x"1b",
x"0f",
x"28",
x"2c",
x"20",
x"3c",
x"39",
x"8d",
x"91",
x"22",
x"11",
x"11",
x"69",
x"9d",
x"a0",
x"a0",
x"a0",
x"a0",
x"b3",
x"cd",
x"d2",
x"5f",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"02",
x"07",
x"0f",
x"20",
x"20",
x"20",
x"20",
x"20",
x"1d",
x"15",
x"2b",
x"2c",
x"20",
x"2a",
x"45",
x"8a",
x"80",
x"17",
x"0b",
x"0b",
x"36",
x"5f",
x"62",
x"62",
x"62",
x"62",
x"82",
x"e2",
x"ff",
x"61",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"0f",
x"20",
x"20",
x"20",
x"20",
x"1c",
x"0e",
x"20",
x"24",
x"23",
x"20",
x"20",
x"45",
x"88",
x"82",
x"20",
x"00",
x"11",
x"1e",
x"27",
x"28",
x"28",
x"28",
x"34",
x"67",
x"dc",
x"ff",
x"61",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"0f",
x"20",
x"20",
x"37",
x"22",
x"1f",
x"1d",
x"20",
x"20",
x"20",
x"20",
x"39",
x"46",
x"88",
x"85",
x"24",
x"00",
x"03",
x"1a",
x"20",
x"20",
x"20",
x"20",
x"22",
x"5c",
x"dc",
x"ff",
x"61",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"0f",
x"20",
x"20",
x"20",
x"39",
x"1f",
x"14",
x"0d",
x"2e",
x"3c",
x"27",
x"39",
x"2a",
x"68",
x"77",
x"20",
x"10",
x"09",
x"16",
x"20",
x"1c",
x"24",
x"32",
x"1e",
x"43",
x"99",
x"ae",
x"53",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"0f",
x"20",
x"20",
x"20",
x"20",
x"1b",
x"02",
x"11",
x"20",
x"20",
x"20",
x"20",
x"3e",
x"37",
x"21",
x"03",
x"03",
x"00",
x"12",
x"33",
x"1e",
x"24",
x"39",
x"32",
x"43",
x"57",
x"3c",
x"10",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"0f",
x"20",
x"20",
x"20",
x"20",
x"1d",
x"11",
x"20",
x"20",
x"20",
x"20",
x"2a",
x"32",
x"1b",
x"08",
x"09",
x"09",
x"08",
x"57",
x"89",
x"95",
x"8b",
x"93",
x"a6",
x"a6",
x"b9",
x"94",
x"3f",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"0f",
x"20",
x"20",
x"20",
x"20",
x"20",
x"20",
x"20",
x"20",
x"20",
x"20",
x"3c",
x"21",
x"20",
x"1b",
x"08",
x"08",
x"1b",
x"54",
x"64",
x"74",
x"73",
x"6d",
x"74",
x"8e",
x"cc",
x"91",
x"24",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"0f",
x"20",
x"20",
x"20",
x"20",
x"23",
x"2e",
x"20",
x"20",
x"20",
x"20",
x"2c",
x"20",
x"20",
x"26",
x"25",
x"1a",
x"20",
x"39",
x"23",
x"22",
x"2d",
x"28",
x"27",
x"48",
x"96",
x"7c",
x"37",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"04",
x"17",
x"20",
x"20",
x"20",
x"21",
x"27",
x"20",
x"20",
x"20",
x"20",
x"20",
x"20",
x"20",
x"2a",
x"32",
x"20",
x"20",
x"27",
x"22",
x"34",
x"20",
x"28",
x"2b",
x"26",
x"3e",
x"76",
x"5b",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"13",
x"20",
x"20",
x"20",
x"20",
x"20",
x"20",
x"20",
x"20",
x"0c",
x"06",
x"06",
x"06",
x"07",
x"09",
x"06",
x"06",
x"1a",
x"20",
x"25",
x"20",
x"22",
x"23",
x"20",
x"20",
x"2e",
x"11",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"01",
x"02",
x"19",
x"1e",
x"1e",
x"1e",
x"1e",
x"10",
x"02",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00"


);

signal car_green: car :=(

x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"05",
x"01",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"0f",
x"03",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"0c",
x"0f",
x"0f",
x"0f",
x"0f",
x"0f",
x"06",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"02",
x"0f",
x"0f",
x"0f",
x"0f",
x"0f",
x"02",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"0d",
x"5b",
x"7d",
x"7e",
x"7e",
x"7e",
x"75",
x"40",
x"09",
x"10",
x"01",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"0c",
x"62",
x"77",
x"75",
x"7e",
x"71",
x"31",
x"02",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"20",
x"36",
x"24",
x"76",
x"a7",
x"a9",
x"a9",
x"a9",
x"99",
x"5c",
x"32",
x"5c",
x"5b",
x"5a",
x"5a",
x"5a",
x"5a",
x"5a",
x"36",
x"05",
x"25",
x"8a",
x"9d",
x"8e",
x"ae",
x"d8",
x"93",
x"2e",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"09",
x"54",
x"82",
x"28",
x"29",
x"36",
x"3b",
x"4a",
x"37",
x"34",
x"2a",
x"4d",
x"a8",
x"b5",
x"b5",
x"b5",
x"b5",
x"b5",
x"b5",
x"6d",
x"21",
x"3d",
x"46",
x"3e",
x"3e",
x"58",
x"b1",
x"a7",
x"5a",
x"15",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"06",
x"13",
x"16",
x"3e",
x"44",
x"43",
x"29",
x"2c",
x"42",
x"33",
x"24",
x"15",
x"23",
x"61",
x"4b",
x"2c",
x"28",
x"28",
x"28",
x"28",
x"25",
x"20",
x"24",
x"22",
x"2c",
x"3d",
x"2e",
x"3c",
x"33",
x"0c",
x"02",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"02",
x"42",
x"95",
x"a0",
x"a0",
x"a0",
x"9c",
x"72",
x"40",
x"64",
x"96",
x"a4",
x"a6",
x"9b",
x"54",
x"0b",
x"0c",
x"0c",
x"00",
x"19",
x"21",
x"37",
x"27",
x"2e",
x"1d",
x"1d",
x"22",
x"87",
x"5c",
x"05",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"08",
x"4a",
x"84",
x"7d",
x"7a",
x"7a",
x"7a",
x"65",
x"2d",
x"59",
x"7e",
x"8b",
x"99",
x"7c",
x"7d",
x"54",
x"0b",
x"05",
x"03",
x"12",
x"1f",
x"1f",
x"17",
x"0e",
x"10",
x"0d",
x"20",
x"5b",
x"42",
x"12",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"18",
x"33",
x"26",
x"20",
x"20",
x"1e",
x"0e",
x"05",
x"21",
x"27",
x"20",
x"30",
x"2a",
x"89",
x"86",
x"1d",
x"0b",
x"06",
x"1f",
x"50",
x"52",
x"42",
x"42",
x"4b",
x"4a",
x"42",
x"52",
x"26",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"0f",
x"20",
x"20",
x"20",
x"20",
x"1b",
x"00",
x"06",
x"18",
x"20",
x"20",
x"20",
x"29",
x"8d",
x"8c",
x"12",
x"0a",
x"11",
x"50",
x"9a",
x"a0",
x"a0",
x"a0",
x"a0",
x"aa",
x"c9",
x"d1",
x"5f",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"0f",
x"20",
x"20",
x"20",
x"20",
x"1b",
x"00",
x"08",
x"25",
x"28",
x"20",
x"20",
x"3b",
x"8e",
x"91",
x"12",
x"06",
x"0b",
x"2d",
x"5e",
x"5f",
x"4d",
x"55",
x"62",
x"82",
x"e0",
x"fb",
x"61",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"0f",
x"20",
x"20",
x"20",
x"1f",
x"06",
x"00",
x"03",
x"18",
x"23",
x"20",
x"20",
x"45",
x"8f",
x"93",
x"12",
x"00",
x"00",
x"19",
x"27",
x"27",
x"20",
x"23",
x"28",
x"5d",
x"d9",
x"fb",
x"61",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"0f",
x"20",
x"20",
x"20",
x"20",
x"18",
x"00",
x"00",
x"10",
x"20",
x"20",
x"20",
x"2c",
x"8f",
x"9c",
x"22",
x"00",
x"00",
x"19",
x"20",
x"20",
x"20",
x"20",
x"20",
x"5a",
x"d9",
x"fb",
x"61",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"0f",
x"20",
x"20",
x"20",
x"20",
x"18",
x"00",
x"00",
x"10",
x"20",
x"20",
x"39",
x"2a",
x"68",
x"6d",
x"10",
x"00",
x"00",
x"16",
x"20",
x"1c",
x"1d",
x"14",
x"0e",
x"43",
x"ab",
x"b2",
x"53",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"0b",
x"1d",
x"1b",
x"18",
x"18",
x"00",
x"00",
x"03",
x"14",
x"20",
x"20",
x"19",
x"3e",
x"37",
x"21",
x"00",
x"00",
x"00",
x"12",
x"33",
x"1e",
x"24",
x"30",
x"26",
x"43",
x"57",
x"3c",
x"10",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"13",
x"12",
x"02",
x"00",
x"00",
x"03",
x"14",
x"20",
x"20",
x"20",
x"0e",
x"32",
x"19",
x"00",
x"00",
x"00",
x"08",
x"57",
x"88",
x"8b",
x"8b",
x"93",
x"a6",
x"ad",
x"bb",
x"94",
x"3f",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"07",
x"19",
x"20",
x"12",
x"0f",
x"0f",
x"14",
x"20",
x"18",
x"11",
x"1c",
x"2d",
x"11",
x"11",
x"0a",
x"00",
x"00",
x"16",
x"48",
x"62",
x"66",
x"73",
x"6d",
x"74",
x"99",
x"cf",
x"91",
x"24",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"06",
x"18",
x"20",
x"20",
x"20",
x"20",
x"20",
x"20",
x"19",
x"13",
x"1d",
x"2c",
x"13",
x"16",
x"1c",
x"13",
x"13",
x"1c",
x"20",
x"20",
x"22",
x"2d",
x"28",
x"27",
x"48",
x"96",
x"7c",
x"27",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"13",
x"20",
x"20",
x"20",
x"20",
x"20",
x"20",
x"20",
x"20",
x"20",
x"0c",
x"1f",
x"20",
x"27",
x"2d",
x"13",
x"19",
x"20",
x"20",
x"20",
x"20",
x"28",
x"2b",
x"26",
x"3e",
x"76",
x"53",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"13",
x"20",
x"20",
x"20",
x"20",
x"20",
x"20",
x"20",
x"10",
x"06",
x"01",
x"05",
x"06",
x"07",
x"09",
x"02",
x"04",
x"1a",
x"20",
x"20",
x"20",
x"22",
x"23",
x"20",
x"20",
x"2e",
x"11",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"01",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"01",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"02",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00"

);

signal car_blue: car :=(


x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"0b",
x"02",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"1e",
x"06",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"18",
x"1e",
x"1e",
x"1e",
x"1e",
x"1e",
x"0b",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"04",
x"1e",
x"1e",
x"1e",
x"1e",
x"1e",
x"05",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"1a",
x"6b",
x"8a",
x"8b",
x"8b",
x"8b",
x"8b",
x"4c",
x"09",
x"20",
x"01",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"0e",
x"6f",
x"8b",
x"8b",
x"8b",
x"80",
x"33",
x"02",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"2a",
x"40",
x"3a",
x"7d",
x"aa",
x"ac",
x"ac",
x"ac",
x"a0",
x"5f",
x"32",
x"64",
x"5b",
x"5a",
x"5a",
x"5a",
x"5a",
x"5a",
x"36",
x"05",
x"39",
x"8b",
x"a3",
x"a9",
x"c0",
x"d3",
x"94",
x"2e",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"12",
x"66",
x"86",
x"50",
x"49",
x"51",
x"52",
x"52",
x"52",
x"4e",
x"44",
x"68",
x"ac",
x"b5",
x"b5",
x"b5",
x"b5",
x"b5",
x"b5",
x"82",
x"3b",
x"42",
x"4d",
x"4f",
x"51",
x"77",
x"b7",
x"bd",
x"74",
x"2b",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"0d",
x"26",
x"25",
x"4a",
x"48",
x"75",
x"4b",
x"48",
x"46",
x"42",
x"44",
x"24",
x"3c",
x"7f",
x"50",
x"4a",
x"45",
x"48",
x"45",
x"44",
x"44",
x"40",
x"40",
x"40",
x"55",
x"78",
x"58",
x"46",
x"4c",
x"11",
x"03",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"04",
x"45",
x"9a",
x"b9",
x"c0",
x"c0",
x"c0",
x"ae",
x"6b",
x"87",
x"c0",
x"c0",
x"c0",
x"ba",
x"6a",
x"24",
x"3b",
x"17",
x"00",
x"33",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"8f",
x"7a",
x"09",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"10",
x"57",
x"92",
x"9a",
x"9a",
x"9a",
x"9a",
x"8e",
x"6d",
x"8e",
x"a1",
x"9a",
x"9a",
x"98",
x"84",
x"78",
x"2c",
x"13",
x"13",
x"28",
x"3e",
x"40",
x"40",
x"40",
x"40",
x"40",
x"32",
x"63",
x"58",
x"25",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"1e",
x"40",
x"40",
x"40",
x"57",
x"40",
x"40",
x"40",
x"61",
x"58",
x"40",
x"40",
x"46",
x"8d",
x"96",
x"40",
x"40",
x"2e",
x"31",
x"64",
x"75",
x"75",
x"75",
x"75",
x"75",
x"5a",
x"6f",
x"34",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"08",
x"22",
x"30",
x"40",
x"40",
x"40",
x"5b",
x"40",
x"40",
x"40",
x"61",
x"58",
x"40",
x"40",
x"46",
x"8d",
x"96",
x"40",
x"40",
x"2c",
x"6c",
x"a1",
x"c0",
x"c0",
x"c0",
x"c0",
x"c0",
x"d8",
x"da",
x"7b",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"05",
x"25",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"61",
x"72",
x"4a",
x"40",
x"6e",
x"b4",
x"ab",
x"2e",
x"17",
x"17",
x"4a",
x"62",
x"6d",
x"6d",
x"6d",
x"6d",
x"86",
x"db",
x"f1",
x"7c",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"16",
x"40",
x"40",
x"40",
x"40",
x"6c",
x"40",
x"40",
x"40",
x"48",
x"4f",
x"44",
x"40",
x"59",
x"ca",
x"b7",
x"39",
x"31",
x"31",
x"3d",
x"40",
x"40",
x"40",
x"40",
x"40",
x"84",
x"df",
x"f0",
x"7c",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"16",
x"40",
x"40",
x"40",
x"6e",
x"7f",
x"70",
x"40",
x"40",
x"5d",
x"78",
x"4e",
x"40",
x"4c",
x"ca",
x"b7",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"6b",
x"d3",
x"f0",
x"7c",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"16",
x"40",
x"40",
x"68",
x"78",
x"78",
x"70",
x"40",
x"40",
x"61",
x"80",
x"7a",
x"78",
x"4e",
x"8a",
x"8c",
x"40",
x"3c",
x"3e",
x"40",
x"40",
x"40",
x"40",
x"40",
x"3c",
x"5f",
x"a1",
x"b1",
x"6c",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"16",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"61",
x"80",
x"50",
x"40",
x"7e",
x"67",
x"40",
x"40",
x"24",
x"30",
x"4c",
x"5d",
x"5c",
x"53",
x"5e",
x"43",
x"44",
x"58",
x"50",
x"11",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"16",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"55",
x"69",
x"4a",
x"40",
x"65",
x"40",
x"40",
x"40",
x"40",
x"40",
x"73",
x"ba",
x"ba",
x"a1",
x"c0",
x"b7",
x"b8",
x"bf",
x"9d",
x"40",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"0c",
x"30",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"5a",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"5b",
x"81",
x"84",
x"84",
x"84",
x"84",
x"a5",
x"d1",
x"ab",
x"26",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"1e",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"57",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"67",
x"a2",
x"88",
x"28",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"1e",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"4b",
x"5a",
x"7b",
x"67",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"05",
x"2a",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"13",
x"10",
x"35",
x"1d",
x"29",
x"29",
x"1d",
x"35",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"4a",
x"17",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"02",
x"2b",
x"3c",
x"3c",
x"3c",
x"3c",
x"3c",
x"3c",
x"3c",
x"3c",
x"08",
x"00",
x"03",
x"01",
x"02",
x"02",
x"01",
x"03",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"04",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00"



);

signal x,y : std_logic_vector (9 downto 0); 
signal redsig: std_logic_vector(7 downto 0);
signal greensig: std_logic_vector(7 downto 0);
signal bluesig: std_logic_vector(7 downto 0);
signal x_decide: std_logic_vector(4 downto 0);
signal y_decide: std_logic_vector(4 downto 0); 
signal calculator, calculator2: std_logic_vector(9 downto 0); 


signal index: std_logic_vector(9 downto 0);
begin



color_process: process(DrawX,DrawY,Car_X_center,Car_Y_center)
begin

x<= DrawX+CONV_STD_LOGIC_VECTOR(20, 10)-Car_X_center;
y<= DrawY+CONV_STD_LOGIC_VECTOR(15, 10)-Car_Y_center;


calculator<= y(4 downto 0) & "00000";
calculator2 <= calculator + (y(6 downto 0) & "000");
index <= calculator2+CONV_STD_LOGIC_VECTOR(39, 10)-x;



-----------------------------------------------------------------------------------
redsig<= car_red(conv_integer(index));		
draw_red<=redsig;    ---Draw the Red parts of the frog if he is moving up
------------------------------------------------------------------------------------
greensig<= car_green(conv_integer( index) );	
draw_green<=greensig;		---Draw the Green parts of the frog if he is moving up. 
----------------------------------------------------------------------------------
bluesig<= car_blue(conv_integer( index));	
draw_blue<=bluesig;		---Draw the blue parts of the frog if he is moving up. 
------------------------------------------------------------------------------------



end process;



end table; 
