library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


entity frog_drawer is 
	Port(
		 
		 DrawX: in std_logic_vector( 9 downto 0); 
		 DrawY: in std_logic_vector( 9 downto 0);
		 Ball_X_center: in std_logic_vector (9 downto 0); 
		 Ball_Y_center: in std_logic_vector (9 downto 0); 
		 keyboard_input : in std_logic_vector(2 downto 0);
		 draw_frog_red: out std_logic_vector(7 downto 0);
		 draw_frog_green: out std_logic_vector(7 downto 0);
		 draw_frog_blue: out std_logic_vector(7 downto 0);
		 frog_life_red: out std_logic_vector(7 downto 0);
		 frog_life_green: out std_logic_vector(7 downto 0);
		 frog_life_blue: out std_logic_vector(7 downto 0)
		 );
end entity;



architecture table of frog_drawer is

type frog is array (1023 downto 0) of std_logic_vector(7 downto 0);
signal red_frog_up : frog := (

x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ab",
x"7c",
x"ca",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"df",
x"5e",
x"76",
x"b9",
x"cf",
x"9c",
x"68",
x"9c",
x"ac",
x"99",
x"7a",
x"f5",
x"ff",
x"ff",
x"ff",
x"ff",
x"c7",
x"5b",
x"a4",
x"ed",
x"ff",
x"ff",
x"ff",
x"ed",
x"5b",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"92",
x"ec",
x"b4",
x"29",
x"00",
x"00",
x"ec",
x"ec",
x"ec",
x"ec",
x"ec",
x"9e",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"ff",
x"ea",
x"58",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"a6",
x"ff",
x"c7",
x"30",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"68",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"77",
x"b7",
x"1c",
x"00",
x"00",
x"ff",
x"ff",
x"dc",
x"86",
x"70",
x"8d",
x"d0",
x"a2",
x"27",
x"00",
x"00",
x"ff",
x"ff",
x"e5",
x"be",
x"ce",
x"62",
x"77",
x"c4",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"9f",
x"c5",
x"10",
x"05",
x"0a",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"df",
x"e2",
x"f3",
x"79",
x"0c",
x"09",
x"97",
x"d8",
x"ef",
x"ff",
x"ff",
x"77",
x"0b",
x"0c",
x"dc",
x"f4",
x"b0",
x"d0",
x"ff",
x"00",
x"00",
x"00",
x"0a",
x"0b",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"f0",
x"f5",
x"ff",
x"78",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"ff",
x"ff",
x"70",
x"00",
x"00",
x"e4",
x"ff",
x"c0",
x"d7",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"eb",
x"eb",
x"f5",
x"65",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"ff",
x"ff",
x"70",
x"00",
x"00",
x"da",
x"f5",
x"b6",
x"d4",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"80",
x"80",
x"50",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"b0",
x"6b",
x"70",
x"1e",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"ff",
x"ff",
x"70",
x"00",
x"00",
x"62",
x"70",
x"50",
x"be",
x"ff",
x"00",
x"00",
x"00",
x"50",
x"80",
x"ff",
x"ff",
x"e1",
x"4d",
x"00",
x"00",
x"ff",
x"ff",
x"80",
x"00",
x"00",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"ff",
x"ff",
x"70",
x"00",
x"00",
x"00",
x"00",
x"00",
x"af",
x"ff",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"ff",
x"e0",
x"4b",
x"00",
x"00",
x"ff",
x"ff",
x"80",
x"00",
x"00",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"ff",
x"ff",
x"70",
x"00",
x"00",
x"00",
x"00",
x"00",
x"af",
x"ff",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"ff",
x"db",
x"46",
x"00",
x"00",
x"1e",
x"ef",
x"7d",
x"0e",
x"0e",
x"0e",
x"0e",
x"36",
x"c7",
x"ff",
x"ff",
x"ff",
x"ff",
x"78",
x"0e",
x"0e",
x"0e",
x"0f",
x"08",
x"a4",
x"ef",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"ff",
x"db",
x"46",
x"00",
x"00",
x"00",
x"00",
x"54",
x"e4",
x"eb",
x"e8",
x"e8",
x"f2",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"f2",
x"e8",
x"e8",
x"e8",
x"ef",
x"80",
x"00",
x"00",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"ff",
x"d1",
x"3a",
x"00",
x"00",
x"00",
x"00",
x"60",
x"eb",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"80",
x"00",
x"00",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"ff",
x"e9",
x"56",
x"00",
x"00",
x"00",
x"00",
x"60",
x"eb",
x"ff",
x"e9",
x"c4",
x"d5",
x"f8",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"8a",
x"06",
x"00",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"ff",
x"ff",
x"e4",
x"cf",
x"cf",
x"cf",
x"cf",
x"c8",
x"eb",
x"ff",
x"42",
x"1e",
x"2f",
x"b9",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"aa",
x"a8",
x"cf",
x"cf",
x"cf",
x"cf",
x"ed",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"e0",
x"eb",
x"ff",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"b0",
x"cd",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"e4",
x"d4",
x"d5",
x"d6",
x"e6",
x"e0",
x"eb",
x"ff",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"b0",
x"cd",
x"da",
x"d5",
x"d4",
x"e4",
x"ff",
x"ff",
x"ff",
x"ff",
x"f6",
x"66",
x"0f",
x"14",
x"17",
x"4e",
x"b0",
x"eb",
x"ff",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"9e",
x"80",
x"26",
x"14",
x"0f",
x"46",
x"db",
x"ff",
x"ff",
x"ff",
x"da",
x"44",
x"00",
x"00",
x"00",
x"00",
x"60",
x"eb",
x"ff",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"80",
x"00",
x"00",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"ff",
x"d8",
x"43",
x"00",
x"00",
x"00",
x"00",
x"60",
x"eb",
x"ff",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"80",
x"00",
x"00",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"ff",
x"db",
x"46",
x"00",
x"00",
x"00",
x"00",
x"33",
x"a7",
x"c4",
x"00",
x"00",
x"00",
x"7a",
x"ac",
x"c4",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"c0",
x"af",
x"62",
x"00",
x"00",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"ff",
x"db",
x"46",
x"00",
x"00",
x"ff",
x"ff",
x"80",
x"00",
x"00",
x"6e",
x"ff",
x"bb",
x"26",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"af",
x"ff",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"ff",
x"e6",
x"53",
x"00",
x"00",
x"ff",
x"ff",
x"80",
x"00",
x"00",
x"88",
x"ff",
x"c7",
x"30",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"af",
x"ff",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"8c",
x"a8",
x"38",
x"00",
x"00",
x"ff",
x"ff",
x"80",
x"00",
x"00",
x"59",
x"dc",
x"a6",
x"2a",
x"00",
x"10",
x"ff",
x"ff",
x"e5",
x"d0",
x"d0",
x"00",
x"00",
x"08",
x"b4",
x"ff",
x"00",
x"00",
x"00",
x"78",
x"8c",
x"50",
x"08",
x"19",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"d7",
x"af",
x"af",
x"0d",
x"3a",
x"29",
x"79",
x"af",
x"b9",
x"ff",
x"ff",
x"8c",
x"32",
x"32",
x"16",
x"af",
x"b4",
x"e9",
x"ff",
x"00",
x"00",
x"00",
x"19",
x"08",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"ff",
x"ff",
x"70",
x"00",
x"00",
x"e3",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"02",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"9d",
x"fb",
x"fb",
x"fb",
x"fa",
x"6d",
x"00",
x"00",
x"7d",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"58",
x"40",
x"2b",
x"04",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"40",
x"40",
x"40",
x"9a",
x"d0",
x"d0",
x"d0",
x"c7",
x"74",
x"40",
x"40",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"28",
x"40",
x"ff",
x"ff",
x"d0",
x"39",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"ff",
x"da",
x"44",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"ff",
x"f4",
x"63",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"31",
x"00",
x"00",
x"9f",
x"ff"


);

signal green_frog_up: frog :=(

x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"cd",
x"ba",
x"e7",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"df",
x"5e",
x"7e",
x"d4",
x"f0",
x"d7",
x"68",
x"9c",
x"ac",
x"99",
x"7a",
x"f5",
x"ff",
x"ff",
x"ff",
x"ff",
x"d7",
x"97",
x"c6",
x"f8",
x"ff",
x"ff",
x"ff",
x"f2",
x"d9",
x"d8",
x"ba",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"92",
x"ec",
x"de",
x"cc",
x"cc",
x"d8",
x"ec",
x"ec",
x"ec",
x"ec",
x"ec",
x"9e",
x"ff",
x"ff",
x"ff",
x"ff",
x"56",
x"e7",
x"c4",
x"e0",
x"ff",
x"ff",
x"ff",
x"ef",
x"e3",
x"ee",
x"d0",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"a6",
x"ff",
x"f1",
x"e0",
x"e0",
x"ee",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"68",
x"ff",
x"ff",
x"ff",
x"ff",
x"6a",
x"fb",
x"d2",
x"e0",
x"ff",
x"ff",
x"9e",
x"d2",
x"ba",
x"e0",
x"c2",
x"ff",
x"ff",
x"d0",
x"5e",
x"40",
x"a5",
x"e8",
x"e4",
x"e0",
x"e0",
x"e0",
x"ff",
x"ff",
x"f2",
x"e8",
x"e8",
x"47",
x"40",
x"a0",
x"ff",
x"ff",
x"6a",
x"f7",
x"cf",
x"e4",
x"c5",
x"4c",
x"d4",
x"c0",
x"cf",
x"e0",
x"c2",
x"ff",
x"ff",
x"84",
x"03",
x"00",
x"8a",
x"f6",
x"e0",
x"f2",
x"e6",
x"fd",
x"ff",
x"ff",
x"ee",
x"e0",
x"fb",
x"38",
x"00",
x"08",
x"b4",
x"ff",
x"6a",
x"f7",
x"df",
x"ce",
x"bf",
x"60",
x"f9",
x"e0",
x"e0",
x"e0",
x"c2",
x"ff",
x"ff",
x"80",
x"00",
x"00",
x"88",
x"f7",
x"e0",
x"f3",
x"ff",
x"ff",
x"ff",
x"ff",
x"ee",
x"e0",
x"e0",
x"35",
x"00",
x"00",
x"af",
x"ff",
x"6a",
x"f7",
x"e0",
x"e0",
x"f9",
x"56",
x"e5",
x"d0",
x"dc",
x"e0",
x"c2",
x"ff",
x"ff",
x"85",
x"11",
x"0b",
x"91",
x"f0",
x"e0",
x"f3",
x"ff",
x"ff",
x"ff",
x"ff",
x"ee",
x"e0",
x"e0",
x"2f",
x"0d",
x"0a",
x"af",
x"ff",
x"6a",
x"f7",
x"e0",
x"d4",
x"e5",
x"a0",
x"dd",
x"b2",
x"b6",
x"e0",
x"c2",
x"ff",
x"ff",
x"b0",
x"81",
x"74",
x"c2",
x"e0",
x"e0",
x"f3",
x"ff",
x"ff",
x"ff",
x"ff",
x"ee",
x"e0",
x"e0",
x"8c",
x"7a",
x"58",
x"b9",
x"ff",
x"6a",
x"f7",
x"d9",
x"d0",
x"dd",
x"ff",
x"ff",
x"e9",
x"d4",
x"e0",
x"c2",
x"ff",
x"ff",
x"db",
x"e1",
x"da",
x"e0",
x"e0",
x"e0",
x"f3",
x"ff",
x"ff",
x"ff",
x"ff",
x"ee",
x"e0",
x"e0",
x"d6",
x"e0",
x"a6",
x"ca",
x"ff",
x"6a",
x"f7",
x"c8",
x"df",
x"ff",
x"ff",
x"ff",
x"ea",
x"d6",
x"e0",
x"c2",
x"ff",
x"ff",
x"d2",
x"d0",
x"e1",
x"e0",
x"e0",
x"e0",
x"f3",
x"ff",
x"ff",
x"ff",
x"ff",
x"ee",
x"e0",
x"e0",
x"e0",
x"ea",
x"a2",
x"c4",
x"ff",
x"50",
x"f7",
x"c4",
x"db",
x"ff",
x"ff",
x"ff",
x"e7",
x"d2",
x"e0",
x"e0",
x"5e",
x"f7",
x"dd",
x"ec",
x"e4",
x"e0",
x"e0",
x"e1",
x"f4",
x"ff",
x"ff",
x"ff",
x"ff",
x"ee",
x"e0",
x"e0",
x"e0",
x"ea",
x"c3",
x"d6",
x"fb",
x"8e",
x"f6",
x"c4",
x"db",
x"ff",
x"ff",
x"ff",
x"e7",
x"d2",
x"e0",
x"e0",
x"c8",
x"c8",
x"d4",
x"f5",
x"eb",
x"e8",
x"e8",
x"f2",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"f2",
x"e8",
x"e8",
x"e8",
x"ef",
x"f4",
x"d2",
x"c8",
x"e0",
x"e0",
x"c4",
x"db",
x"ff",
x"ff",
x"ff",
x"dd",
x"cd",
x"ee",
x"e1",
x"e0",
x"e0",
x"e0",
x"f5",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ea",
x"e0",
x"e0",
x"e4",
x"d2",
x"e0",
x"ff",
x"ff",
x"ff",
x"ed",
x"d4",
x"c9",
x"b9",
x"b8",
x"b8",
x"cc",
x"f5",
x"ff",
x"ec",
x"ec",
x"ec",
x"f8",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ec",
x"c2",
x"b8",
x"b8",
x"c0",
x"bc",
x"d8",
x"ff",
x"ff",
x"ff",
x"ff",
x"f8",
x"ef",
x"ed",
x"ed",
x"ed",
x"da",
x"ed",
x"ff",
x"e0",
x"e0",
x"e0",
x"f3",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"c6",
x"cf",
x"ed",
x"ed",
x"ef",
x"ee",
x"f6",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"e0",
x"eb",
x"ff",
x"e0",
x"e0",
x"e0",
x"f3",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"b0",
x"cd",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"eb",
x"db",
x"e1",
x"e1",
x"ea",
x"e3",
x"ed",
x"ff",
x"e0",
x"e0",
x"e0",
x"f3",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"b3",
x"cf",
x"e5",
x"e1",
x"e0",
x"eb",
x"ff",
x"ff",
x"ff",
x"ff",
x"fa",
x"b0",
x"73",
x"83",
x"84",
x"a2",
x"e3",
x"f5",
x"ff",
x"e0",
x"e0",
x"e0",
x"f3",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"d2",
x"d2",
x"91",
x"84",
x"82",
x"a5",
x"f1",
x"ff",
x"ff",
x"ff",
x"e5",
x"d9",
x"da",
x"d2",
x"d2",
x"d2",
x"d9",
x"f5",
x"ff",
x"e0",
x"e0",
x"e0",
x"f3",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"f8",
x"dc",
x"d2",
x"d2",
x"da",
x"d5",
x"e2",
x"ff",
x"ff",
x"ff",
x"e4",
x"d3",
x"e2",
x"e0",
x"e3",
x"f0",
x"e0",
x"f5",
x"ff",
x"e0",
x"e0",
x"e0",
x"f3",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ea",
x"f4",
x"e0",
x"e2",
x"cc",
x"de",
x"ff",
x"ff",
x"ff",
x"e7",
x"d2",
x"e0",
x"e0",
x"a4",
x"a5",
x"c2",
x"e1",
x"e2",
x"e0",
x"e0",
x"e0",
x"e1",
x"e2",
x"e2",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"e2",
x"e2",
x"d3",
x"ae",
x"a6",
x"c4",
x"e0",
x"c4",
x"db",
x"ff",
x"ff",
x"ff",
x"e7",
x"d2",
x"e0",
x"c2",
x"ff",
x"ff",
x"de",
x"e7",
x"e4",
x"e2",
x"ff",
x"f1",
x"e0",
x"e0",
x"e0",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"e0",
x"ea",
x"b0",
x"cd",
x"ff",
x"6a",
x"f7",
x"c4",
x"db",
x"ff",
x"ff",
x"ff",
x"ef",
x"db",
x"e0",
x"c2",
x"ff",
x"ff",
x"d5",
x"d6",
x"e1",
x"e2",
x"ff",
x"f1",
x"e0",
x"e0",
x"e0",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"e8",
x"ea",
x"b0",
x"cd",
x"ff",
x"6a",
x"f7",
x"c4",
x"db",
x"ff",
x"ff",
x"a9",
x"c4",
x"cb",
x"e0",
x"c2",
x"ff",
x"ff",
x"d0",
x"c1",
x"b4",
x"e1",
x"f0",
x"e9",
x"e0",
x"e0",
x"e0",
x"ff",
x"ff",
x"f7",
x"f0",
x"f0",
x"dc",
x"ca",
x"a0",
x"cd",
x"ff",
x"6a",
x"f7",
x"cb",
x"c4",
x"a9",
x"92",
x"b0",
x"b7",
x"cf",
x"e0",
x"c2",
x"ff",
x"ff",
x"eb",
x"de",
x"d9",
x"a4",
x"f0",
x"e0",
x"ed",
x"f5",
x"f5",
x"ff",
x"ff",
x"ee",
x"e0",
x"e0",
x"77",
x"e4",
x"dc",
x"ef",
x"ff",
x"6a",
x"f7",
x"dc",
x"c2",
x"b0",
x"60",
x"f5",
x"de",
x"e0",
x"e0",
x"c2",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"88",
x"f7",
x"e0",
x"f3",
x"ff",
x"ff",
x"ff",
x"ff",
x"ee",
x"e0",
x"e0",
x"ea",
x"ff",
x"ff",
x"ff",
x"ff",
x"6a",
x"f7",
x"e0",
x"de",
x"f5",
x"60",
x"fb",
x"ee",
x"de",
x"e0",
x"c2",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"a2",
x"f2",
x"e9",
x"fa",
x"fb",
x"fb",
x"fb",
x"fb",
x"fa",
x"f9",
x"f9",
x"97",
x"ff",
x"ff",
x"ff",
x"ff",
x"6a",
x"f7",
x"e0",
x"ef",
x"f9",
x"88",
x"cb",
x"a6",
x"ba",
x"e0",
x"c2",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"8b",
x"b8",
x"b8",
x"c7",
x"d0",
x"d0",
x"d0",
x"d0",
x"c2",
x"b8",
x"b8",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"6a",
x"f7",
x"d9",
x"c1",
x"b8",
x"ff",
x"ff",
x"d7",
x"bf",
x"e0",
x"c2",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"6a",
x"f7",
x"c4",
x"db",
x"ff",
x"ff",
x"ff",
x"e1",
x"d6",
x"f3",
x"d6",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"6a",
x"fc",
x"d7",
x"e3",
x"ff",
x"ff",
x"ff",
x"f6",
x"c9",
x"b2",
x"94",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"65",
x"b2",
x"a1",
x"d4",
x"ff"

);

signal blue_frog_up: frog :=(

x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ab",
x"8f",
x"c1",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"c2",
x"00",
x"2e",
x"a1",
x"c3",
x"9c",
x"14",
x"68",
x"68",
x"41",
x"03",
x"f5",
x"ff",
x"ff",
x"ff",
x"ff",
x"c9",
x"6f",
x"a6",
x"ed",
x"ff",
x"ff",
x"ff",
x"ed",
x"5b",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"89",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"ff",
x"ea",
x"58",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"40",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"64",
x"b7",
x"1c",
x"00",
x"00",
x"ff",
x"ff",
x"d0",
x"7f",
x"70",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"46",
x"70",
x"b8",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"9f",
x"c8",
x"10",
x"03",
x"0a",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"de",
x"e2",
x"f3",
x"38",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"c0",
x"f3",
x"a0",
x"c7",
x"ff",
x"00",
x"00",
x"00",
x"0a",
x"0b",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"e0",
x"eb",
x"ff",
x"78",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"c8",
x"ff",
x"c0",
x"d7",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"d6",
x"d7",
x"eb",
x"65",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"b4",
x"eb",
x"ac",
x"d1",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"80",
x"80",
x"50",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"a0",
x"56",
x"60",
x"1e",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"44",
x"60",
x"40",
x"b9",
x"ff",
x"00",
x"00",
x"00",
x"50",
x"80",
x"ff",
x"ff",
x"e1",
x"4d",
x"00",
x"00",
x"ff",
x"ff",
x"80",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"af",
x"ff",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"ff",
x"ea",
x"58",
x"00",
x"00",
x"ff",
x"ff",
x"80",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"af",
x"ff",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"ff",
x"e7",
x"54",
x"00",
x"00",
x"1c",
x"e1",
x"71",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"a4",
x"ef",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"ff",
x"e7",
x"54",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"ff",
x"dd",
x"48",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"ff",
x"ed",
x"5b",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"ff",
x"ff",
x"e4",
x"cf",
x"cf",
x"cf",
x"cf",
x"68",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"8e",
x"cf",
x"cf",
x"cf",
x"cf",
x"ed",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"80",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"af",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"e4",
x"cf",
x"cf",
x"d1",
x"e6",
x"7f",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"af",
x"d5",
x"cf",
x"cf",
x"e3",
x"fe",
x"ff",
x"ff",
x"ff",
x"f6",
x"66",
x"00",
x"00",
x"05",
x"4a",
x"4b",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"6d",
x"14",
x"00",
x"00",
x"42",
x"d7",
x"ff",
x"ff",
x"ff",
x"da",
x"44",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"ff",
x"e1",
x"4d",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"ff",
x"e7",
x"54",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"ff",
x"e7",
x"54",
x"00",
x"00",
x"ff",
x"ff",
x"80",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"af",
x"ff",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"ff",
x"ef",
x"5d",
x"00",
x"00",
x"ff",
x"ff",
x"80",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"af",
x"ff",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"8c",
x"a8",
x"38",
x"00",
x"00",
x"ff",
x"ff",
x"80",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"af",
x"ff",
x"00",
x"00",
x"00",
x"78",
x"8c",
x"50",
x"08",
x"19",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"d7",
x"af",
x"af",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"16",
x"af",
x"af",
x"e6",
x"ff",
x"00",
x"00",
x"00",
x"19",
x"08",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"e3",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"00",
x"97",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"00",
x"00",
x"40",
x"40",
x"28",
x"00",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"40",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"28",
x"40",
x"ff",
x"ff",
x"c9",
x"31",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"ff",
x"e1",
x"4d",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"00",
x"00",
x"00",
x"9f",
x"ff",
x"ff",
x"ff",
x"f6",
x"66",
x"00",
x"00",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"ff",
x"31",
x"00",
x"00",
x"9f",
x"ff"



);

signal x,y : std_logic_vector (9 downto 0); 
signal redsig: std_logic_vector(7 downto 0);
signal greensig: std_logic_vector(7 downto 0);
signal bluesig: std_logic_vector(7 downto 0);
signal x_decide: std_logic_vector(4 downto 0);
signal y_decide: std_logic_vector(4 downto 0); 


signal index, index2: std_logic_vector(9 downto 0);
signal keyboard_prev: std_logic_vector(1 downto 0); 
begin



color_process: process(DrawX,DrawY,Ball_X_center,Ball_Y_center, keyboard_input)
begin

x<= DrawX+CONV_STD_LOGIC_VECTOR(16, 10)-Ball_X_center;
y<= DrawY+CONV_STD_LOGIC_VECTOR(16, 10)-Ball_Y_center;

x_decide <= x(4 downto 0);
y_decide <= y(4 downto 0); 

if(keyboard_input= "100") then			--Last key pressed was a W
keyboard_prev<= "00";
elsif(keyboard_input= "101") then 		--Last Key pressed was an S
keyboard_prev<= "01";
elsif(keyboard_input= "110") then		--Last Key pressed was an A
keyboard_prev<="10";
elsif(keyboard_input= "111") then		--Last Key pressed was a D
keyboard_prev<="11"; 
end if; 


if(keyboard_prev= "00") then
index<= (not(y_decide)+'1') & x_decide;					--Up


elsif(keyboard_prev= "01") then
index<= y_decide & x_decide;							--Down


elsif(keyboard_prev= "10") then
index<= (not(x_decide)+'1') & y_decide;		--Left    


elsif(keyboard_prev= "11") then
index<= x_decide & y_decide; 							--Right
end if; 
--index<= x_decide & y_decide;
-----------------------------------------------------------------------------------
redsig<= red_frog_up(conv_integer(index));		
draw_frog_red<=redsig;    ---Draw the Red parts of the frog if he is moving up
------------------------------------------------------------------------------------
greensig<= green_frog_up(conv_integer( index) );	
draw_frog_green<=greensig;		---Draw the Green parts of the frog if he is moving up. 
----------------------------------------------------------------------------------
bluesig<= blue_frog_up(conv_integer( index));	
draw_frog_blue<=bluesig;		---Draw the blue parts of the frog if he is moving up. 
------------------------------------------------------------------------------------

index2<= (not(y_decide)+'1') & x_decide;

-----------------------------------------------------------------------------------
frog_life_red<= red_frog_up(conv_integer(index));		
draw_frog_red<=redsig;    ---Draw the Red parts of the frog if he is moving up
------------------------------------------------------------------------------------
frog_life_green<= green_frog_up(conv_integer( index) );	
draw_frog_green<=greensig;		---Draw the Green parts of the frog if he is moving up. 
----------------------------------------------------------------------------------
frog_life_blue<= blue_frog_up(conv_integer( index));	
draw_frog_blue<=bluesig;		---Draw the blue parts of the frog if he is moving up. 
------------------------------------------------------------------------------------



end process;



end table; 
