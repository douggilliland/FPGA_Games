module	spi	(
			input	MOSI,
			input	clk,
			input	SS,
			output	MISO
		);
endmodule
