library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package Images is

	-- Tipo das imagens das tiles
	type image_array_t is array(15 downto 0, 15 downto 0) of unsigned(11 downto 0);
	
	-- Imagem de uma caixa
	constant tile_box : image_array_t := (
		(X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0"),
		(X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0"),
		(X"fb0",X"fb0",X"960",X"960",X"960",X"960",X"960",X"960",X"960",X"960",X"960",X"960",X"960",X"960",X"fb0",X"fb0"),
		(X"fb0",X"fb0",X"960",X"960",X"960",X"960",X"960",X"960",X"960",X"960",X"960",X"fb0",X"fb0",X"960",X"fb0",X"fb0"),
		(X"fb0",X"fb0",X"960",X"960",X"960",X"960",X"960",X"960",X"960",X"960",X"fb0",X"fb0",X"fb0",X"960",X"fb0",X"fb0"),
		(X"fb0",X"fb0",X"960",X"960",X"960",X"960",X"960",X"960",X"960",X"fb0",X"fb0",X"fb0",X"960",X"960",X"fb0",X"fb0"),
		(X"fb0",X"fb0",X"960",X"960",X"960",X"960",X"960",X"960",X"fb0",X"fb0",X"fb0",X"960",X"960",X"960",X"fb0",X"fb0"),
		(X"fb0",X"fb0",X"960",X"960",X"960",X"960",X"960",X"fb0",X"fb0",X"fb0",X"960",X"960",X"960",X"960",X"fb0",X"fb0"),
		(X"fb0",X"fb0",X"960",X"960",X"960",X"960",X"fb0",X"fb0",X"fb0",X"960",X"960",X"960",X"960",X"960",X"fb0",X"fb0"),
		(X"fb0",X"fb0",X"960",X"960",X"960",X"fb0",X"fb0",X"fb0",X"960",X"960",X"960",X"960",X"960",X"960",X"fb0",X"fb0"),
		(X"fb0",X"fb0",X"960",X"960",X"fb0",X"fb0",X"fb0",X"960",X"960",X"960",X"960",X"960",X"960",X"960",X"fb0",X"fb0"),
		(X"fb0",X"fb0",X"960",X"fb0",X"fb0",X"fb0",X"960",X"960",X"960",X"960",X"960",X"960",X"960",X"960",X"fb0",X"fb0"),
		(X"fb0",X"fb0",X"960",X"fb0",X"fb0",X"960",X"960",X"960",X"960",X"960",X"960",X"960",X"960",X"960",X"fb0",X"fb0"),
		(X"fb0",X"fb0",X"960",X"960",X"960",X"960",X"960",X"960",X"960",X"960",X"960",X"960",X"960",X"960",X"fb0",X"fb0"),
		(X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0"),
		(X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0",X"fb0")
	);

	-- Imagem de uma caixa sobre um objetivo
	constant tile_box_objective : image_array_t := (
		(X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0"),
		(X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0"),
		(X"dc0",X"dc0",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"dc0",X"dc0"),
		(X"dc0",X"dc0",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"dc0",X"dc0",X"ab1",X"dc0",X"dc0"),
		(X"dc0",X"dc0",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"dc0",X"dc0",X"dc0",X"ab1",X"dc0",X"dc0"),
		(X"dc0",X"dc0",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"dc0",X"dc0",X"dc0",X"ab1",X"ab1",X"dc0",X"dc0"),
		(X"dc0",X"dc0",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"dc0",X"dc0",X"dc0",X"ab1",X"ab1",X"ab1",X"dc0",X"dc0"),
		(X"dc0",X"dc0",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"dc0",X"dc0",X"dc0",X"ab1",X"ab1",X"ab1",X"ab1",X"dc0",X"dc0"),
		(X"dc0",X"dc0",X"ab1",X"ab1",X"ab1",X"ab1",X"dc0",X"dc0",X"dc0",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"dc0",X"dc0"),
		(X"dc0",X"dc0",X"ab1",X"ab1",X"ab1",X"dc0",X"dc0",X"dc0",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"dc0",X"dc0"),
		(X"dc0",X"dc0",X"ab1",X"ab1",X"dc0",X"dc0",X"dc0",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"dc0",X"dc0"),
		(X"dc0",X"dc0",X"ab1",X"dc0",X"dc0",X"dc0",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"dc0",X"dc0"),
		(X"dc0",X"dc0",X"ab1",X"dc0",X"dc0",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"dc0",X"dc0"),
		(X"dc0",X"dc0",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"ab1",X"dc0",X"dc0"),
		(X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0"),
		(X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0",X"dc0")
	);

	-- Imagem do chão
	constant tile_floor : image_array_t := (
		(X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb"),
		(X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb"),
		(X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb"),
		(X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb"),
		(X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb"),
		(X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb"),
		(X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb"),
		(X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb"),
		(X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb"),
		(X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb"),
		(X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb"),
		(X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb"),
		(X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb"),
		(X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb"),
		(X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb"),
		(X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb")
	);

	-- Imagem do objetivo
	constant tile_objective : image_array_t := (
		(X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb"),
		(X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb"),
		(X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb"),
		(X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb"),
		(X"ba7",X"dcb",X"dcb",X"dcb",X"2b4",X"2b4",X"2b4",X"2b4",X"2b4",X"2b4",X"2b4",X"2b4",X"ba7",X"dcb",X"dcb",X"dcb"),
		(X"ba7",X"dcb",X"dcb",X"dcb",X"2b4",X"2b4",X"2b4",X"2b4",X"2b4",X"2b4",X"2b4",X"2b4",X"ba7",X"dcb",X"dcb",X"dcb"),
		(X"ba7",X"dcb",X"dcb",X"dcb",X"2b4",X"2b4",X"2b4",X"2b4",X"2b4",X"2b4",X"2b4",X"2b4",X"ba7",X"dcb",X"dcb",X"dcb"),
		(X"ba7",X"dcb",X"dcb",X"dcb",X"2b4",X"2b4",X"2b4",X"2b4",X"2b4",X"2b4",X"2b4",X"2b4",X"ba7",X"dcb",X"dcb",X"dcb"),
		(X"ba7",X"dcb",X"dcb",X"dcb",X"2b4",X"2b4",X"2b4",X"2b4",X"2b4",X"2b4",X"2b4",X"2b4",X"ba7",X"dcb",X"dcb",X"dcb"),
		(X"ba7",X"dcb",X"dcb",X"dcb",X"2b4",X"2b4",X"2b4",X"2b4",X"2b4",X"2b4",X"2b4",X"2b4",X"ba7",X"dcb",X"dcb",X"dcb"),
		(X"ba7",X"dcb",X"dcb",X"dcb",X"2b4",X"2b4",X"2b4",X"2b4",X"2b4",X"2b4",X"2b4",X"2b4",X"ba7",X"dcb",X"dcb",X"dcb"),
		(X"ba7",X"dcb",X"dcb",X"dcb",X"2b4",X"2b4",X"2b4",X"2b4",X"2b4",X"2b4",X"2b4",X"2b4",X"ba7",X"dcb",X"dcb",X"dcb"),
		(X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb"),
		(X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb"),
		(X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb"),
		(X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb")
	);

	-- Imagem do player
	constant tile_player : image_array_t := (
		(X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb"),
		(X"ba7",X"666",X"666",X"666",X"666",X"666",X"666",X"666",X"666",X"666",X"666",X"666",X"666",X"666",X"666",X"dcb"),
		(X"ba7",X"666",X"666",X"666",X"666",X"666",X"666",X"666",X"666",X"666",X"666",X"666",X"666",X"666",X"666",X"dcb"),
		(X"ba7",X"666",X"666",X"333",X"333",X"333",X"333",X"333",X"333",X"333",X"333",X"333",X"333",X"666",X"666",X"dcb"),
		(X"ba7",X"666",X"666",X"333",X"333",X"333",X"333",X"333",X"333",X"333",X"333",X"333",X"333",X"666",X"666",X"dcb"),
		(X"ba7",X"666",X"666",X"333",X"333",X"333",X"333",X"333",X"333",X"333",X"333",X"333",X"333",X"666",X"666",X"dcb"),
		(X"ba7",X"666",X"666",X"333",X"333",X"333",X"333",X"e12",X"e12",X"333",X"333",X"333",X"333",X"666",X"666",X"dcb"),
		(X"ba7",X"666",X"666",X"333",X"333",X"333",X"e12",X"e12",X"e12",X"e12",X"333",X"333",X"333",X"666",X"666",X"dcb"),
		(X"ba7",X"666",X"666",X"333",X"333",X"333",X"e12",X"e12",X"e12",X"e12",X"333",X"333",X"333",X"666",X"666",X"dcb"),
		(X"ba7",X"666",X"666",X"333",X"333",X"333",X"333",X"e12",X"e12",X"333",X"333",X"333",X"333",X"666",X"666",X"dcb"),
		(X"ba7",X"666",X"666",X"333",X"333",X"333",X"333",X"333",X"333",X"333",X"333",X"333",X"333",X"666",X"666",X"dcb"),
		(X"ba7",X"666",X"666",X"333",X"333",X"333",X"333",X"333",X"333",X"333",X"333",X"333",X"333",X"666",X"666",X"dcb"),
		(X"ba7",X"666",X"666",X"333",X"333",X"333",X"333",X"333",X"333",X"333",X"333",X"333",X"333",X"666",X"666",X"dcb"),
		(X"ba7",X"666",X"666",X"666",X"666",X"666",X"666",X"666",X"666",X"666",X"666",X"666",X"666",X"666",X"666",X"dcb"),
		(X"ba7",X"666",X"666",X"666",X"666",X"666",X"666",X"666",X"666",X"666",X"666",X"666",X"666",X"666",X"666",X"dcb"),
		(X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb",X"ba7",X"dcb",X"dcb",X"dcb")
	);

	-- Imagem de uma parede
	constant tile_wall : image_array_t := (
		(X"fff",X"fff",X"fff",X"fff",X"fff",X"fff",X"fff",X"777",X"fff",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"777"),
		(X"fff",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"777",X"fff",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"777"),
		(X"fff",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"777",X"fff",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"777"),
		(X"fff",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"777",X"fff",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"777"),
		(X"fff",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"777",X"fff",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"777"),
		(X"fff",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"777",X"fff",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"777"),
		(X"fff",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"777",X"fff",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"777"),
		(X"fff",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"777",X"777",X"777",X"777",X"777",X"777",X"777",X"777",X"777"),
		(X"fff",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"777",X"fff",X"fff",X"fff",X"fff",X"fff",X"fff",X"fff",X"777"),
		(X"fff",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"777",X"fff",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"777"),
		(X"fff",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"777",X"fff",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"777"),
		(X"fff",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"777",X"fff",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"777"),
		(X"fff",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"777",X"fff",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"777"),
		(X"fff",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"777",X"fff",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"777"),
		(X"fff",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"777",X"fff",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"777"),
		(X"777",X"777",X"777",X"777",X"777",X"777",X"777",X"777",X"fff",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"ccc",X"777")
	);

	-- Imagem de um check (simbolo de vitória)
	constant check_img : image_array_t := (
		(X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000"),
		(X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000"),
		(X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"9f5",X"000",X"000",X"000",X"000",X"000",X"000",X"000"),
		(X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"9f5",X"000",X"000",X"000",X"000",X"000",X"000"),
		(X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"9f5",X"000",X"000",X"000",X"000",X"000"),
		(X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"9f5",X"9f5",X"000",X"000",X"000",X"000"),
		(X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"9f5",X"9f5",X"9f5",X"000",X"000",X"000"),
		(X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"9f5",X"9f5",X"9f5",X"000",X"000",X"000",X"000"),
		(X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"9f5",X"9f5",X"9f5",X"000",X"000",X"000",X"000",X"000"),
		(X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"9f5",X"9f5",X"9f5",X"000",X"000",X"000",X"000",X"000",X"000"),
		(X"000",X"000",X"000",X"000",X"000",X"000",X"9f5",X"9f5",X"9f5",X"000",X"000",X"000",X"000",X"000",X"000",X"000"),
		(X"000",X"000",X"000",X"000",X"000",X"9f5",X"9f5",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000"),
		(X"000",X"000",X"000",X"000",X"9f5",X"9f5",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000"),
		(X"000",X"000",X"000",X"9f5",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000"),
		(X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000"),
		(X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000",X"000")
	);

end package;
