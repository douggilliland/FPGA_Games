module microfono
(
	input             CLK,
	input      	  D_IN,
	output            BCLK,
	output            WS,
	output            SELECT,
	output            DONE,
	output     [17:0] D_OUT,

);
endmodule
