----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 26.01.2017 10:52:07
-- Design Name: 
-- Module Name: CellArray - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library work; 
use work.TableType.ALL;

entity CellArray is
    Generic ( HEIGHT : integer := 60;
              WIDTH : integer := 80);
    Port ( CLK : in STD_LOGIC;
           CLK_SLOW : in STD_LOGIC;
           RST : in STD_LOGIC;
           STATE : out TABLE(WIDTH downto 1, HEIGHT downto 1));
end CellArray;

architecture Behavioral of CellArray is

signal tableNumber : integer range 0 to 4 := 0;

--constant voidTable : TABLE(33 downto 0, 25 downto 0)  := ((others=> (others=>'0')));
--constant voidTable : TABLE(41 downto 0, 31 downto 0)  := ((others=> (others=>'0')));
--constant voidTable : TABLE(65 downto 0, 49 downto 0)  := ((others=> (others=>'0')));

--constant initTable : TABLE(33 downto 0, 25 downto 0)  := 
--   ("00000000000000000000000000",
--    "00100000000000000000000000",
--    "00010000000000000000000000",
--    "01110000000000000000000000",
--    "00000000000000000000000000",
--    "00000000000000000000000000",
--    "00000000000000000000000000",
--    "00000000000000000000000000",
--    "00000000000000000000000000",
--    "00000000000000000000000000",
--    "00000000000000000000000000",
--    "00000000000000000000000000",
--    "00000000000000000000000000",
--    "00000000000000000000000000",
--    "00000000000000000000000000",
--    "00000000000000000000000000",
--    "00000000000000000000000000",
--    "00000000000000000000000000",
--    "00000000000000000000000000",
--    "00000000000000000000000000",
--    "00000000000000000000000000",
--    "00000000000000000000000000",
--    "00000000000000000000000000",
--    "00000000000000000000000000",
--    "00000000000000000000000000",
--    "00000000000000000000000000",
--    "00000000000000000000000000",
--    "00000000000000000000000000",
--    "00000000000000000000000000",
--    "00000000000000000000000000",
--    "00000000000000000000000000",
--    "00000000000000000000000000",
--    "00000000000000000000000000",
--    "00000000000000000000000000");
--constant initTable : TABLE(41 downto 0, 31 downto 0)  := 
--    ("00000000000000000000000000000000",
--     "00000000000000000000000000000000",
--     "00000000000000000000000011000000",
--     "00000000000000000000000011000000",
--     "00000000000000000000000000000000",
--     "00000000000000000000000000000000",
--     "00000000000000000000000000000000",
--     "00000000000000000000000000000000",
--     "00000000000000000000000000000000",
--     "00000000000000000000000000000000",
--     "00000000000000000000000000000000",
--     "00000000000000000000000000000000",
--     "00000000000000000000000111000000",
--     "00000000000000000000001000100000",
--     "00000000000000000000010000010000",
--     "00000000000000000000010000010000",
--     "00000000000000000000000010000000",
--     "00000000000000000000001000100000",
--     "00000000000000000000000111000000",
--     "00000000000000000000000010000000",
--     "00000000000000000000000000000000",
--     "00000000000000000000000000000000",
--     "00000000000000000000000001110000",
--     "00000000000000000000000001110000",
--     "00000000000000000000000010001000",
--     "00000000000000000000000000000000",
--     "00000000000000000000000110001100",
--     "00000000000000000000000000000000",
--     "00000000000000000000000000000000",
--     "00000000000000000000000000000000",
--     "00000000000000000000000000000000",
--     "00000000000000000000000000000000",
--     "00000000000000000000000000000000",
--     "00000000000000000000000000000000",
--     "00000000000000000000000000000000",
--     "00000000000000000000000000000000",
--     "00000000000000000000000000110000",
--     "00000000000000000000000000110000",
--     "00000000000000000000000000000000",
--     "00000000000000000000000000000000",
--     "00000000000000000000000000000000",
--     "00000000000000000000000000000000");
--constant initTable : TABLE(65 downto 0, 49 downto 0)  := 
--   ("00000000000000000000000000000000000000000000000000",
--    "00100000000000000000000000000000000000000000000000",
--    "00010000000000000000000000000000000000000000000000",
--    "01110000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000");
signal initTable : TABLE(81 downto 0, 61 downto 0)  := 
   ("00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00010000000000000000000000000000000000000000000000000000000000",
    "00001000000000000000000000000000000000000000000000000000000000",
    "00111000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000");
    

constant initTable0 : TABLE(81 downto 0, 61 downto 0)  := 
   ("00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00010000000000000000000000000000000000000000000000000000000000",
    "00001000000000000000000000000000000000000000000000000000000000",
    "00111000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000");

constant initTable1 : TABLE(81 downto 0, 61 downto 0)  := 
   ("00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000100000000000000000000000000000",
    "00000000000000000000000000000000101000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000010000000000000000000000000000",
    "00000000000000000000000000000000100000000000000000000000000000",
    "00000000000000000000000000000000100000000000000000000000000000",
    "00000000000000000000000000000000100000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000");


constant initTable2 : TABLE(81 downto 0, 61 downto 0)  := 
   ("00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000011000000000000000000000000000",
    "00000000000000000000000000000000110000000000000000000000000000",
    "00000000000000000000000000000000010000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000");


constant initTable3 : TABLE(81 downto 0, 61 downto 0)  := 
    ("00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000011000000",
     "00000000000000000000000000000000000000000000000000000011000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000111000000",
     "00000000000000000000000000000000000000000000000000001000100000",
     "00000000000000000000000000000000000000000000000000010000010000",
     "00000000000000000000000000000000000000000000000000010000010000",
     "00000000000000000000000000000000000000000000000000000010000000",
     "00000000000000000000000000000000000000000000000000001000100000",
     "00000000000000000000000000000000000000000000000000000111000000",
     "00000000000000000000000000000000000000000000000000000010000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000001110000",
     "00000000000000000000000000000000000000000000000000000001110000",
     "00000000000000000000000000000000000000000000000000000010001000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000110001100",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000110000",
     "00000000000000000000000000000000000000000000000000000000110000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000",
     "00000000000000000000000000000000000000000000000000000000000000");


constant initTable4 : TABLE(81 downto 0, 61 downto 0)  := 
   ("00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00010000000000000000000000000000000000000000000000000000000000",
    "00001000000000000000000000000000000000000000000000000000000000",
    "00111000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000000000000000000");



--constant initTable : TABLE(129 downto 0, 97 downto 0)  := 
--   ("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "01110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
--    "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");
    
signal internalState : TABLE(WIDTH+1 downto 0, HEIGHT+1 downto 0) := initTable;

component Cell is
    generic (CELL_INIT : STD_LOGIC := '0');
    Port ( CLK : in STD_LOGIC;
           CLK_E : in STD_LOGIC;
           PROX : in STD_LOGIC_VECTOR(7 downto 0);
           RST : in STD_LOGIC;
           RST_VALUE : in STD_LOGIC;
           STATE : out STD_LOGIC);
end component;
 
begin

-- Using a generate loop for the Cell matrix
MAPGEN: FOR i IN 1 TO WIDTH generate
    LINGEN: FOR j IN 1 TO HEIGHT generate
         CellX : Cell generic map (initTable1(i,j)) port map (CLK => CLK,      
                                                 CLK_E => CLK_SLOW,
                                                 PROX => (internalState(i+1,j)&internalState(i+1,j+1)&internalState(i,j+1)&internalState(i-1,j+1)&internalState(i-1,j)&internalState(i-1,j-1)&internalState(i,j-1)&internalState(i+1,j-1)),
                                                 RST => RST,
                                                 RST_VALUE => initTable(i,j),
                                                 STATE => internalState(i,j));
    end generate LINGEN;
end generate MAPGEN;

-- Connect internalState to STATE output. FOR LOOP needs to be in a process. 
process(internalState)
begin
STATE_CONNECT_LINE: FOR i IN 1 TO WIDTH loop
    STATE_CONNECT_CELL: FOR j IN 1 TO HEIGHT loop
        STATE(i,j) <= internalState(i,j);
    end loop STATE_CONNECT_CELL;
end loop STATE_CONNECT_LINE;
end process;

process(RST) -- reset button changes the original map between 5 maps
begin
if (RST = '1' AND RST'EVENT) then
    if (tableNumber = 0) then 
        initTable <= initTable1;
        tableNumber <= tableNumber+1;
    elsif (tableNumber = 1) then
        initTable <= initTable1;
        tableNumber <= tableNumber+1;
    elsif (tableNumber = 2) then
        initTable <= initTable2;
        tableNumber <= tableNumber+1;
    elsif (tableNumber = 3) then
        initTable <= initTable3;
        tableNumber <= tableNumber+1;
    elsif (tableNumber = 4) then
        initTable <= initTable4;
        tableNumber <= 0;
    end if;
end if;
end process;

end Behavioral;
