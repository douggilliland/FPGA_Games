module contador		(
				output wire	[7:0] count,
				output reg	calculate,
				input	ECHO,
				input	CLKOUT,
				input	reset
			);
	reg [7:0] count0;
	reg logico;
	//reg calculate;
	initial 
	begin
		count0=0;
		//pulse=0;
		calculate=0;
	end
	
	always@(posedge CLKOUT)
	begin
		logico=(count0[7]||count0[6]||count0[5]||count0[4]||count0[3]||count0[2]||count0[1]||count0[0]);
		if(reset)
		begin
			count0=0;
			calculate=0;
		end
		else
		begin
			//	Cuenta el rango que tiene el pulso del ECHO del sensor
			//
			if(ECHO)
			begin
				count0=count0+1;
			end
			if(!ECHO && logico)
			begin
				calculate = 1;
			end
		end
	end
	assign count = count0;
endmodule
