----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    10:13:59 05/25/2015 
-- Design Name: 
-- Module Name:    SCORE_ROM - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity SCORE_ROM is
 Port ( Hposition   : in  STD_LOGIC_VECTOR(10 downto 0);
		  Vposition   : in  STD_LOGIC_VECTOR(9 downto 0);
		  VIDON       : in  STD_LOGIC;
		  enable_game : in  STD_LOGIC;
        obj_rgb     : out  STD_LOGIC;
		  obj_on      : out  STD_LOGIC );
end SCORE_ROM;

architecture Behavioral of SCORE_ROM is

type ROM is array(0 to 39) of std_logic_vector(99 downto 0);
constant content : ROM := (

0 =>"1111111111111111110000111111111111111100001111111111111100001111111111111000000011111111111111111100",
1 =>"1111111111111111110001111111111111111100011111111111111110001111111111111100000011111111111111111100",
2 =>"1111111111111111110011111111111111111100111111111111111111001111111111111110000011111111111111111100",
3 =>"1111111111111111110011111111000000000000111111111111111111001111111111111110000011111100000000000000",
4 =>"1111110000000000000011111110000000000000111110000000111111001111110000111111000011111100000000000000",
5 =>"1111110000000000000011111110000000000000111110000000011111001111110000111111000011111100000000000000",
6 =>"1111110000000000000011111110000000000000111110000000011111001111110000011111100011111100000000000000",
7 =>"1111110000000000000011111110000000000000111110000000011111000111111000011111100011111100000000000000",
8 =>"1111110000000000000011111110000000000000111110000000011111001111110000001111110011111100000000000000",
9 =>"0111111000000000000011111110000000000000111110000000011111001111110000001111110011111100000000000000",
10=>"0011111100000000000011111110000000000000111110000000011111001111110000001111110011111100000000000000",
11=>"0001111110000000000011111110000000000000111110000000011111001111110000001111110011111100000000000000",
12=>"0000111111000000000011111110000000000000111110000000011111001111110000001111110011111100000000000000",
13=>"0000111111000000000011111110000000000000111110000000011111001111110000011111100011111100000000000000",
14=>"0000011111100000000011111110000000000000111110000000011111001111110000111111000011111100000000000000",
15=>"0000011111100000000011111110000000000000111110000000011111001111110000111111100011111100000000000000",
16=>"0000001111110000000011111110000000000000111110000000011111001111111111111110000011111100000000000000",
17=>"0000001111110000000011111110000000000000111110000000011111001111111111111100000011111100000000000000",
18=>"0000000111111000000001111110000000000000111110000000011111001111111111111000000011111100000000000000",
19=>"0000000111111000000011111110000000000000111110000000011111001111111111110000000011111111111110000000",
20=>"0000000011111100000011111110000000000000111110000000011111001111111111100000000011111111111110000000",
21=>"0000000011111100000011111110000000000000111110000000011111001111111111110000000011111111111110000000",
22=>"0000000001111110000011111110000000000000111110000000011111001111110111111000000011111100000000000000",
23=>"0000000001111110000011111110000000000000111110000000011111001111110111111000000011111100000000000000",
24=>"0000000001111110000011111110000000000000111110000000011111001111110011111100000011111100000000000000",
25=>"0000000000111111000011111110000000000000111110000000011111001111110011111100000011111100000000000000",
26=>"0000000000011111100011111110000000000000111110000000011111001111110001111110000011111100000000000000",
27=>"0000000000011111100011111110000000000000111110000000011111001111110001111110000011111100000000000000",
28=>"0000000000001111110011111110000000000000111110000000011111001111110000111111000011111100000000000000",
29=>"0000000000001111110011111110000000000000111110000000011111001111110000011111100011111100000000000000",
30=>"0000000000001111110011111110000000000000111110000000011111001111110000001111110011111100000000000000",
31=>"0000000000001111110011111110000000000000111110000000011111001111110000001111110011111100000000000000",
32=>"0000000000001111110011111110000000000000111110000000011111001111110000001111110011111100000000000000",
33=>"0000000000001111110011111110000000000000111110000000011111001111110000001111110011111100000000000000",
34=>"0000000000001111110011111110000000000000111110000000011111001111110000001111110011111100000000000000",
35=>"0000000000001111110011111110000000000000111110000000011111001111110000001111110011111100000000000000",
36=>"0000000000001111110011111111000000000000111111000000111111001111110000001111110011111111111111111100",
37=>"1111111111111111110011111111111111111100111111111111111111001111110000001111110011111111111111111100",
38=>"1111111111111111110001111111111111111100011111111111111110001111110000001111110011111111111111111100",
39=>"1111111111111111110000111111111111111100001111111111111100001111110000001111110011111111111111111100"
);

signal data_line : std_logic_vector(0 to 99);

constant Hstart : std_logic_vector(10 downto 0) := "01000111111"; -- 575
constant Hend :std_logic_vector(10 downto 0)    := "01010100011"; -- 675
constant Vstart : std_logic_vector(9 downto 0)  := "0000110010"; -- 50
constant Vend : std_logic_vector(9 downto 0)    := "0001011010"; -- 90

signal obj_row :  STD_LOGIC_VECTOR (10 downto 0);
signal obj_col :  STD_LOGIC_VECTOR (9 downto 0);

signal obj_on_sig : std_logic := '0';
signal object_rgb : std_logic := '0';

begin

process(VIDON, enable_game, Hposition, Vposition)

begin

    object_rgb <= '0';
	 obj_on_sig <='0';
	 
	 if VIDON = '1' and enable_game = '1' then
	     
		  	  if (Hposition >= Hstart and Hposition < Hend) and 
	           (Vposition >= Vstart and Vposition < Vend) then
		  
					  obj_on_sig <= '1';
					  obj_row <= (Hposition-Hstart);
					  obj_col <= (Vposition-Vstart);
					  
					  data_line <= content(conv_integer(obj_col));
		  
		           object_rgb <= data_line(conv_integer(obj_row));
					  
		     end if;
		  
	 end if;

end process;
obj_rgb <= object_rgb;
obj_on <= obj_on_sig;

end Behavioral;
